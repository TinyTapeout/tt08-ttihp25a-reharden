* NGSPICE file created from core_prel_parax.ext - technology: sky130A

.subckt core_prel_parax VDD Vbgr VSS
X0 w_18582_n15452.t12 Vbgr.t5 VSS.t52 w_18582_n15452.t11 sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=10
X1 a_19776_n11398# a_20010_n12050# VSS.t30 sky130_fd_pr__res_xhigh_po_0p69 l=1.26
X2 VDD.t33 w_18582_n15452.t13 MINUS.t3 VDD.t32 sky130_fd_pr__pfet_01v8_lvt ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X3 VDD.t56 VDD.t53 VDD.t55 VDD.t54 sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=10
X4 VDD.t52 VDD.t49 VDD.t51 VDD.t50 sky130_fd_pr__pfet_01v8_lvt ad=1.45 pd=10.58 as=0 ps=0 w=5 l=0.5
X5 VSS.t69 VSS.t100 XQ2[0|0].Emitter sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X6 VSS.t72 VSS.t99 XQ2[0|0].Emitter sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X7 VSS.t57 VSS.t98 XQ2[0|0].Emitter sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X8 VSS.t54 VSS.t97 XQ2[0|0].Emitter sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X9 a_19776_n11398# a_19542_n12050# VSS.t40 sky130_fd_pr__res_xhigh_po_0p69 l=1.26
X10 a_12755_n6044# PLUS.t5 VSS.t39 sky130_fd_pr__res_xhigh_po_0p35 l=1
X11 Sop Gcm2 VSS.t15 VSS.t14 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.5
X12 a_13419_n6044# a_13087_n6644# VSS.t41 sky130_fd_pr__res_xhigh_po_0p35 l=1
X13 VSS.t8 VSS.t9 VSS.t7 sky130_fd_pr__res_xhigh_po_0p69 l=1.26
X14 Vbgr.t3 w_18582_n15452.t14 VDD.t31 VDD.t30 sky130_fd_pr__pfet_01v8_lvt ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X15 a_12921_n6044# a_13253_n6644# VSS.t16 sky130_fd_pr__res_xhigh_po_0p35 l=1
X16 w_18582_n15452.t4 Gcm1.t6 VDD.t58 VDD.t57 sky130_fd_pr__pfet_01v8_lvt ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X17 VDD.t48 VDD.t45 VDD.t47 VDD.t46 sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=10
X18 w_18582_n15452.t10 Vbgr.t6 VSS.t49 w_18582_n15452.t9 sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=10
X19 VSS.t13 Gcm2 Sop VSS.t12 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.5
X20 a_13419_n6044# a_13914_n6644# VSS.t3 sky130_fd_pr__res_xhigh_po_0p35 l=1
X21 VSS.t72 VSS.t96 XQ2[0|0].Emitter sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X22 VSS.t60 VSS.t95 XQ2[0|0].Emitter sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X23 VDD.t29 w_18582_n15452.t15 Gcm2 VDD.t28 sky130_fd_pr__pfet_01v8_lvt ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X24 w_18582_n15452.t8 Vbgr.t7 VSS.t50 w_18582_n15452.t7 sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=10
X25 MINUS.t0 a_14080_n6644# VSS.t25 sky130_fd_pr__res_xhigh_po_0p35 l=1
X26 VSS.t94 VSS.t92 Sop VSS.t93 sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.58 as=1.16 ps=8.29 w=8 l=4
X27 VSS.t46 VSS.t47 VSS.t45 sky130_fd_pr__res_xhigh_po_0p35 l=1.05
X28 MINUS.t2 w_18582_n15452.t16 VDD.t27 VDD.t26 sky130_fd_pr__pfet_01v8_lvt ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X29 w_18582_n15452.t6 Vbgr.t8 VSS.t51 w_18582_n15452.t5 sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=10
X30 VDD.t25 w_18582_n15452.t17 MINUS.t1 VDD.t24 sky130_fd_pr__pfet_01v8_lvt ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X31 a_19308_n11398# a_19074_n12050# VSS.t28 sky130_fd_pr__res_xhigh_po_0p69 l=1.26
X32 VDD.t23 w_18582_n15452.t18 Vbgr.t2 VDD.t22 sky130_fd_pr__pfet_01v8_lvt ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X33 Sop VSS.t89 VSS.t91 VSS.t90 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.29 as=2.32 ps=16.58 w=8 l=4
X34 VSS.t69 VSS.t88 XQ2[0|0].Emitter sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X35 VSS.t24 a_12589_n6644# VSS.t23 sky130_fd_pr__res_xhigh_po_0p35 l=1
X36 VSS.t57 VSS.t87 XQ2[0|0].Emitter sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X37 VSS.t69 VSS.t86 XQ2[0|0].Emitter sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X38 Gcm2 w_18582_n15452.t19 VDD.t21 VDD.t20 sky130_fd_pr__pfet_01v8_lvt ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X39 PLUS.t4 w_18582_n15452.t20 VDD.t19 VDD.t18 sky130_fd_pr__pfet_01v8_lvt ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X40 VSS.t54 VSS.t85 XQ2[0|0].Emitter sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X41 a_19308_n11398# a_19542_n12050# VSS.t18 sky130_fd_pr__res_xhigh_po_0p69 l=1.26
X42 Sop PLUS.t6 Gcm1.t5 VSS.t31 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=4
X43 a_12755_n6044# a_13087_n6644# VSS.t105 sky130_fd_pr__res_xhigh_po_0p35 l=1
X44 VDD.t44 VDD.t42 VDD.t44 VDD.t43 sky130_fd_pr__pfet_01v8_lvt ad=0.725 pd=5.29 as=0 ps=0 w=5 l=0.5
X45 MINUS.t4 w_18582_n15452.t21 VDD.t17 VDD.t16 sky130_fd_pr__pfet_01v8_lvt ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X46 VSS.t69 VSS.t84 XQ2[0|0].Emitter sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X47 Vbgr.t4 a_20478_n12050# VSS.t104 sky130_fd_pr__res_xhigh_po_0p69 l=1.26
X48 a_13748_n6044# a_13253_n6644# VSS.t5 sky130_fd_pr__res_xhigh_po_0p35 l=1
X49 VSS.t102 VSS.t103 VSS.t101 sky130_fd_pr__res_xhigh_po_0p35 l=1.05
X50 VDD.t41 VDD.t39 w_18582_n15452.t1 VDD.t40 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=0.58 ps=4.29 w=4 l=1
X51 VSS.t57 VSS.t83 XQ2[0|0].Emitter sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X52 VSS.t60 VSS.t82 XQ2[0|0].Emitter sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X53 VSS.t60 VSS.t81 XQ2[0|0].Emitter sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X54 VSS.t54 VSS.t80 XQ2[0|0].Emitter sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X55 VDD.t15 w_18582_n15452.t22 PLUS.t3 VDD.t14 sky130_fd_pr__pfet_01v8_lvt ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X56 PLUS.t0 XQ2[0|0].Emitter VSS.t4 sky130_fd_pr__res_xhigh_po_0p35 l=1.05
X57 a_14246_n6044# a_13914_n6644# VSS.t44 sky130_fd_pr__res_xhigh_po_0p35 l=1
X58 VSS.t72 VSS.t79 XQ2[0|0].Emitter sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X59 a_13748_n6044# a_14080_n6644# VSS.t43 sky130_fd_pr__res_xhigh_po_0p35 l=1
X60 a_20244_n11398# a_20478_n12050# VSS.t0 sky130_fd_pr__res_xhigh_po_0p69 l=1.26
X61 w_18582_n15452.t3 VDD.t36 VDD.t38 VDD.t37 sky130_fd_pr__pfet_01v8_lvt ad=0.58 pd=4.29 as=1.16 ps=8.58 w=4 l=1
X62 VSS.t60 VSS.t78 XQ2[0|0].Emitter sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X63 Vbgr.t1 w_18582_n15452.t23 VDD.t13 VDD.t12 sky130_fd_pr__pfet_01v8_lvt ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X64 VSS.t2 a_18606_n12050# VSS.t1 sky130_fd_pr__res_xhigh_po_0p69 l=1.26
X65 Sop MINUS.t6 w_18582_n15452.t0 VSS.t17 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=4
X66 VSS.t20 VSS.t21 VSS.t19 sky130_fd_pr__res_xhigh_po_0p35 l=1
X67 VDD.t11 w_18582_n15452.t24 PLUS.t2 VDD.t10 sky130_fd_pr__pfet_01v8_lvt ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X68 a_18840_n11398# a_18606_n12050# VSS.t35 sky130_fd_pr__res_xhigh_po_0p69 l=1.26
X69 PLUS.t1 w_18582_n15452.t25 VDD.t9 VDD.t8 sky130_fd_pr__pfet_01v8_lvt ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X70 VSS.t69 VSS.t77 XQ2[0|0].Emitter sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X71 VSS.t33 VSS.t34 VSS.t32 sky130_fd_pr__res_xhigh_po_0p35 l=1
X72 VDD.t7 w_18582_n15452.t26 Vbgr.t0 VDD.t6 sky130_fd_pr__pfet_01v8_lvt ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X73 VSS.t72 VSS.t76 XQ2[0|0].Emitter sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X74 VSS.t57 VSS.t75 XQ2[0|0].Emitter sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X75 VSS.t54 VSS.t74 XQ2[0|0].Emitter sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X76 VSS.t72 VSS.t73 XQ2[0|0].Emitter sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X77 a_18840_n11398# a_19074_n12050# VSS.t22 sky130_fd_pr__res_xhigh_po_0p69 l=1.26
X78 Gcm1.t3 Gcm1.t2 VDD.t60 VDD.t59 sky130_fd_pr__pfet_01v8_lvt ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X79 Gcm1.t4 PLUS.t7 Sop VSS.t42 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=4
X80 a_20244_n11398# a_20010_n12050# VSS.t48 sky130_fd_pr__res_xhigh_po_0p69 l=1.26
X81 VSS.t69 VSS.t68 MINUS.t5 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X82 VDD.t5 w_18582_n15452.t27 Gcm2 VDD.t4 sky130_fd_pr__pfet_01v8_lvt ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X83 VDD.t35 Gcm1.t7 w_18582_n15452.t2 VDD.t34 sky130_fd_pr__pfet_01v8_lvt ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X84 VSS.t72 VSS.t71 XQ2[0|0].Emitter sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X85 VSS.t60 VSS.t70 XQ2[0|0].Emitter sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X86 Gcm2 Gcm2 VSS.t11 VSS.t10 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.5
X87 VSS.t67 VSS.t64 VSS.t66 VSS.t65 sky130_fd_pr__nfet_01v8_lvt ad=0.58 pd=4.58 as=0 ps=0 w=2 l=0.5
X88 a_12921_n6044# a_12589_n6644# VSS.t6 sky130_fd_pr__res_xhigh_po_0p35 l=1
X89 VSS.t63 VSS.t61 Gcm2 VSS.t62 sky130_fd_pr__nfet_01v8_lvt ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.5
X90 a_14246_n6044# VSS.t27 VSS.t26 sky130_fd_pr__res_xhigh_po_0p35 l=1
X91 VSS.t60 VSS.t59 XQ2[0|0].Emitter sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X92 VDD.t1 Gcm1.t0 Gcm1.t1 VDD.t0 sky130_fd_pr__pfet_01v8_lvt ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X93 VSS.t37 VSS.t38 VSS.t36 sky130_fd_pr__res_xhigh_po_0p69 l=1.26
X94 Gcm2 w_18582_n15452.t28 VDD.t3 VDD.t2 sky130_fd_pr__pfet_01v8_lvt ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X95 VSS.t57 VSS.t58 XQ2[0|0].Emitter sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X96 VSS.t57 VSS.t56 XQ2[0|0].Emitter sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X97 VSS.t54 VSS.t55 XQ2[0|0].Emitter sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X98 VSS.t54 VSS.t53 XQ2[0|0].Emitter sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X99 w_18582_n15452.t0 MINUS.t7 Sop VSS.t29 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=4
R0 Vbgr.n3 Vbgr.n1 166.519
R1 Vbgr.n3 Vbgr.n2 166.518
R2 Vbgr Vbgr.t4 21.9643
R3 Vbgr.n2 Vbgr.t0 5.7135
R4 Vbgr.n2 Vbgr.t3 5.7135
R5 Vbgr.n1 Vbgr.t2 5.7135
R6 Vbgr.n1 Vbgr.t1 5.7135
R7 Vbgr.n7 Vbgr.t6 4.97522
R8 Vbgr.n9 Vbgr.t5 4.9198
R9 Vbgr.n8 Vbgr.t8 4.9198
R10 Vbgr.n7 Vbgr.t7 4.9198
R11 Vbgr.n10 Vbgr.n9 4.63261
R12 Vbgr.n6 Vbgr.n5 2.75531
R13 Vbgr.n5 Vbgr.n3 2.24383
R14 Vbgr.n5 Vbgr.n4 0.994731
R15 Vbgr.n11 Vbgr 0.871594
R16 Vbgr.n11 Vbgr.n10 0.391125
R17 Vbgr.n6 Vbgr 0.253909
R18 Vbgr Vbgr.n0 0.245692
R19 Vbgr.n4 Vbgr 0.143857
R20 Vbgr.n10 Vbgr.n6 0.114136
R21 Vbgr.n6 Vbgr.n0 0.0774231
R22 Vbgr.n9 Vbgr.n8 0.0559149
R23 Vbgr.n8 Vbgr.n7 0.0559149
R24 Vbgr.n4 Vbgr.n0 0.0293462
R25 Vbgr Vbgr.n11 0.0197308
R26 VSS.n341 VSS.n340 727100
R27 VSS.n1185 VSS.n3 78819
R28 VSS.n5287 VSS.n341 38374.9
R29 VSS.n5285 VSS.n344 36926.8
R30 VSS.n1182 VSS.n1169 12208.2
R31 VSS.n5503 VSS.n58 10933.5
R32 VSS.n5286 VSS.n5285 8231.18
R33 VSS.n5287 VSS.n5286 8171.97
R34 VSS.n5283 VSS.n344 7702.65
R35 VSS.n5282 VSS.n347 5618.46
R36 VSS.n4013 VSS.n1162 5394.32
R37 VSS.n5284 VSS.n5283 4019.23
R38 VSS.n5288 VSS.n339 3874.21
R39 VSS.n5510 VSS.n48 3091.12
R40 VSS.n1188 VSS.n48 3091.12
R41 VSS.n1188 VSS.n1186 3091.12
R42 VSS.n5285 VSS.n5284 3088.46
R43 VSS.n1184 VSS.n344 3008.04
R44 VSS.n5288 VSS.n5287 2988.68
R45 VSS.n1184 VSS.n1183 1829.32
R46 VSS.n5282 VSS.n5281 1818.78
R47 VSS.n5510 VSS.n47 1814.52
R48 VSS.n945 VSS.n944 1801.72
R49 VSS.n2996 VSS.n2995 1801.72
R50 VSS.n2817 VSS.n2816 1801.72
R51 VSS.n2929 VSS.n2928 1801.72
R52 VSS.n944 VSS.n903 1559.06
R53 VSS.n912 VSS.n903 1559.06
R54 VSS.n913 VSS.n912 1559.06
R55 VSS.n930 VSS.n929 1559.06
R56 VSS.n929 VSS.n842 1559.06
R57 VSS.n4546 VSS.n842 1559.06
R58 VSS.n4547 VSS.n4546 1559.06
R59 VSS.n4548 VSS.n4547 1559.06
R60 VSS.n3035 VSS.n2996 1559.06
R61 VSS.n3035 VSS.n3034 1559.06
R62 VSS.n3034 VSS.n3033 1559.06
R63 VSS.n3002 VSS.n3001 1559.06
R64 VSS.n3002 VSS.n1461 1559.06
R65 VSS.n3051 VSS.n1461 1559.06
R66 VSS.n3052 VSS.n3051 1559.06
R67 VSS.n3053 VSS.n3052 1559.06
R68 VSS.n2842 VSS.n2817 1559.06
R69 VSS.n2842 VSS.n2841 1559.06
R70 VSS.n2841 VSS.n2840 1559.06
R71 VSS.n3113 VSS.n1427 1559.06
R72 VSS.n3114 VSS.n3113 1559.06
R73 VSS.n3117 VSS.n3114 1559.06
R74 VSS.n3117 VSS.n3116 1559.06
R75 VSS.n3116 VSS.n3115 1559.06
R76 VSS.n2961 VSS.n2929 1559.06
R77 VSS.n2961 VSS.n2960 1559.06
R78 VSS.n2960 VSS.n2959 1559.06
R79 VSS.n2930 VSS.n1445 1559.06
R80 VSS.n3080 VSS.n1445 1559.06
R81 VSS.n3081 VSS.n3080 1559.06
R82 VSS.n3083 VSS.n3081 1559.06
R83 VSS.n3083 VSS.n3082 1559.06
R84 VSS.n1180 VSS.n1179 1286.03
R85 VSS.n1186 VSS.n47 1276.61
R86 VSS.n1172 VSS.n1170 1257.25
R87 VSS.n4395 VSS.n963 1135.73
R88 VSS.n1524 VSS.n247 1135.73
R89 VSS.n2527 VSS.n343 1135.73
R90 VSS.n4327 VSS.n963 1105.64
R91 VSS.n5290 VSS.n247 1105.64
R92 VSS.n2288 VSS.n345 1105.64
R93 VSS.n5286 VSS.n343 1090.6
R94 VSS.n5069 VSS.n5068 1083.5
R95 VSS.n3997 VSS.n3996 854.934
R96 VSS.n5284 VSS.n345 834.872
R97 VSS.n1186 VSS.n1185 829.258
R98 VSS.n930 VSS.t69 814.173
R99 VSS.n3001 VSS.t69 814.173
R100 VSS.n1427 VSS.t69 814.173
R101 VSS.n2930 VSS.t69 814.173
R102 VSS.n913 VSS.t69 744.883
R103 VSS.n3033 VSS.t69 744.883
R104 VSS.n2840 VSS.t69 744.883
R105 VSS.n2959 VSS.t69 744.883
R106 VSS.n4071 VSS.n4 676.923
R107 VSS.n4099 VSS.n4071 676.923
R108 VSS.n4099 VSS.n4098 676.923
R109 VSS.n4098 VSS.n4097 676.923
R110 VSS.n4097 VSS.n4072 676.923
R111 VSS.n4088 VSS.n4087 676.923
R112 VSS.n4087 VSS.n4086 676.923
R113 VSS.n4326 VSS.n4325 676.923
R114 VSS.n4327 VSS.n4326 676.923
R115 VSS.n4395 VSS.n4394 676.923
R116 VSS.n4394 VSS.n4393 676.923
R117 VSS.n4393 VSS.n4334 676.923
R118 VSS.n4362 VSS.n4334 676.923
R119 VSS.n4362 VSS.n4361 676.923
R120 VSS.n4351 VSS.n4350 676.923
R121 VSS.n4351 VSS.n338 676.923
R122 VSS.n5291 VSS.n5289 676.923
R123 VSS.n5291 VSS.n5290 676.923
R124 VSS.n1525 VSS.n1524 676.923
R125 VSS.n2558 VSS.n1525 676.923
R126 VSS.n2558 VSS.n2557 676.923
R127 VSS.n2557 VSS.n2556 676.923
R128 VSS.n2556 VSS.n1526 676.923
R129 VSS.n2547 VSS.n2546 676.923
R130 VSS.n2546 VSS.n2545 676.923
R131 VSS.n2545 VSS.n1535 676.923
R132 VSS.n2536 VSS.n1535 676.923
R133 VSS.n2536 VSS.n342 676.923
R134 VSS.n2527 VSS.n2526 676.923
R135 VSS.n2526 VSS.n2525 676.923
R136 VSS.n2525 VSS.n1564 676.923
R137 VSS.n2234 VSS.n1564 676.923
R138 VSS.n2234 VSS.n2233 676.923
R139 VSS.n2246 VSS.n2245 676.923
R140 VSS.n2246 VSS.n2224 676.923
R141 VSS.n2286 VSS.n2224 676.923
R142 VSS.n2287 VSS.n2286 676.923
R143 VSS.n2288 VSS.n2287 676.923
R144 VSS.n2297 VSS.n346 676.923
R145 VSS.n2297 VSS.n2126 676.923
R146 VSS.n2310 VSS.n2126 676.923
R147 VSS.n2311 VSS.n2310 676.923
R148 VSS.n2312 VSS.n2311 676.923
R149 VSS.n2314 VSS.n2119 676.923
R150 VSS.n2327 VSS.n2119 676.923
R151 VSS.n2328 VSS.n2327 676.923
R152 VSS.n2329 VSS.n2328 676.923
R153 VSS.n2329 VSS.n347 676.923
R154 VSS.n57 VSS.n52 640.297
R155 VSS.n5504 VSS.n52 637.191
R156 VSS.n5505 VSS.n51 635.47
R157 VSS.n4325 VSS.n3 631.795
R158 VSS.n56 VSS.n51 627.563
R159 VSS.n1168 VSS.n3 585.779
R160 VSS.n4144 VSS.n45 585
R161 VSS.n4145 VSS.n4144 585
R162 VSS.n4144 VSS.n61 585
R163 VSS.n5262 VSS.n5261 585
R164 VSS.n5261 VSS.n5260 585
R165 VSS.n5263 VSS.n359 585
R166 VSS.n359 VSS.n358 585
R167 VSS.n5265 VSS.n5264 585
R168 VSS.n5266 VSS.n5265 585
R169 VSS.n357 VSS.n356 585
R170 VSS.n5267 VSS.n357 585
R171 VSS.n5270 VSS.n5269 585
R172 VSS.n5269 VSS.n5268 585
R173 VSS.n5271 VSS.n354 585
R174 VSS.n354 VSS.n353 585
R175 VSS.n5273 VSS.n5272 585
R176 VSS.n5274 VSS.n5273 585
R177 VSS.n355 VSS.n351 585
R178 VSS.n5275 VSS.n351 585
R179 VSS.n5277 VSS.n352 585
R180 VSS.n5277 VSS.n5276 585
R181 VSS.n5278 VSS.n348 585
R182 VSS.n5281 VSS.n5280 585
R183 VSS.n4982 VSS.n4953 585
R184 VSS.n4986 VSS.n4953 585
R185 VSS.n4984 VSS.n4983 585
R186 VSS.n4985 VSS.n4984 585
R187 VSS.n4981 VSS.n4956 585
R188 VSS.n4956 VSS.n4955 585
R189 VSS.n4980 VSS.n4979 585
R190 VSS.n4979 VSS.n4978 585
R191 VSS.n4976 VSS.n4957 585
R192 VSS.n4977 VSS.n4976 585
R193 VSS.n4975 VSS.n4959 585
R194 VSS.n4975 VSS.n4974 585
R195 VSS.n4969 VSS.n4958 585
R196 VSS.n4973 VSS.n4958 585
R197 VSS.n4971 VSS.n4970 585
R198 VSS.n4972 VSS.n4971 585
R199 VSS.n4968 VSS.n4961 585
R200 VSS.n4961 VSS.n4960 585
R201 VSS.n612 VSS.n608 585
R202 VSS.n5010 VSS.n612 585
R203 VSS.n5008 VSS.n5007 585
R204 VSS.n5009 VSS.n5008 585
R205 VSS.n5006 VSS.n617 585
R206 VSS.n617 VSS.n616 585
R207 VSS.n5005 VSS.n5004 585
R208 VSS.n5004 VSS.n5003 585
R209 VSS.n619 VSS.n618 585
R210 VSS.n5002 VSS.n619 585
R211 VSS.n5000 VSS.n4999 585
R212 VSS.n5001 VSS.n5000 585
R213 VSS.n4998 VSS.n623 585
R214 VSS.n623 VSS.n622 585
R215 VSS.n4997 VSS.n4996 585
R216 VSS.n4996 VSS.n4995 585
R217 VSS.n625 VSS.n624 585
R218 VSS.n4994 VSS.n625 585
R219 VSS.n2293 VSS.n674 585
R220 VSS.n2294 VSS.n2221 585
R221 VSS.n2221 VSS.n710 585
R222 VSS.n2294 VSS.n2293 585
R223 VSS.n2293 VSS.n710 585
R224 VSS.n378 VSS.n377 585
R225 VSS.n5236 VSS.n378 585
R226 VSS.n5239 VSS.n5238 585
R227 VSS.n5238 VSS.n5237 585
R228 VSS.n5240 VSS.n376 585
R229 VSS.n376 VSS.n375 585
R230 VSS.n5242 VSS.n5241 585
R231 VSS.n5243 VSS.n5242 585
R232 VSS.n372 VSS.n371 585
R233 VSS.n5244 VSS.n372 585
R234 VSS.n5247 VSS.n5246 585
R235 VSS.n5246 VSS.n5245 585
R236 VSS.n5248 VSS.n369 585
R237 VSS.n369 VSS.n368 585
R238 VSS.n5250 VSS.n5249 585
R239 VSS.n5251 VSS.n5250 585
R240 VSS.n370 VSS.n366 585
R241 VSS.n5252 VSS.n366 585
R242 VSS.n5230 VSS.n381 585
R243 VSS.n5230 VSS.n383 585
R244 VSS.n5230 VSS.n5229 585
R245 VSS.n4967 VSS.n4966 585
R246 VSS.n4966 VSS.n4965 585
R247 VSS.n4963 VSS.n4962 585
R248 VSS.n4964 VSS.n4963 585
R249 VSS.n5232 VSS.n5231 585
R250 VSS.n5231 VSS.n379 585
R251 VSS.n5234 VSS.n5233 585
R252 VSS.n5235 VSS.n5234 585
R253 VSS.n2926 VSS.n2621 585
R254 VSS.n2926 VSS.n2925 585
R255 VSS.n404 VSS.n402 585
R256 VSS.n5223 VSS.n404 585
R257 VSS.n1926 VSS.n674 585
R258 VSS.n2175 VSS.n710 585
R259 VSS.n5228 VSS.n391 585
R260 VSS.n5228 VSS.n5227 585
R261 VSS.n5229 VSS.n5228 585
R262 VSS.n5226 VSS.n391 585
R263 VSS.n5227 VSS.n5226 585
R264 VSS.n5226 VSS.n5225 585
R265 VSS.n5224 VSS.n402 585
R266 VSS.n5224 VSS.n5223 585
R267 VSS.n5225 VSS.n5224 585
R268 VSS.n3224 VSS.n1345 585
R269 VSS.n3256 VSS.n3224 585
R270 VSS.n3224 VSS.n3223 585
R271 VSS.n4554 VSS.n838 585
R272 VSS.n4555 VSS.n4554 585
R273 VSS.n4554 VSS.n4550 585
R274 VSS.n4549 VSS.n838 585
R275 VSS.n4550 VSS.n4549 585
R276 VSS.n946 VSS.n900 585
R277 VSS.n4407 VSS.n946 585
R278 VSS.n949 VSS.n244 585
R279 VSS.n3254 VSS.n244 585
R280 VSS.n2923 VSS.n244 585
R281 VSS.n251 VSS.n244 585
R282 VSS.n5372 VSS.n266 585
R283 VSS.n5372 VSS.n279 585
R284 VSS.n5372 VSS.n285 585
R285 VSS.n1521 VSS.n290 585
R286 VSS.n5372 VSS.n290 585
R287 VSS.n1521 VSS.n251 585
R288 VSS.n5372 VSS.n251 585
R289 VSS.n4470 VSS.n406 585
R290 VSS.n5221 VSS.n406 585
R291 VSS.n2530 VSS.n406 585
R292 VSS.n3188 VSS.n407 585
R293 VSS.n1623 VSS.n407 585
R294 VSS.n2531 VSS.n1561 585
R295 VSS.n1561 VSS.n407 585
R296 VSS.n2531 VSS.n2530 585
R297 VSS.n2530 VSS.n407 585
R298 VSS.n3222 VSS.n1355 585
R299 VSS.n3222 VSS.n3221 585
R300 VSS.n3223 VSS.n3222 585
R301 VSS.n3215 VSS.n406 585
R302 VSS.n1387 VSS.n406 585
R303 VSS.n3220 VSS.n1355 585
R304 VSS.n3221 VSS.n3220 585
R305 VSS.n3220 VSS.n456 585
R306 VSS.n3217 VSS.n454 585
R307 VSS.n3218 VSS.n456 585
R308 VSS.n5120 VSS.n503 585
R309 VSS.n606 VSS.n605 585
R310 VSS.n614 VSS.n613 585
R311 VSS.n5014 VSS.n610 585
R312 VSS.n5011 VSS.n610 585
R313 VSS.n5014 VSS.n5013 585
R314 VSS.n5013 VSS.n5012 585
R315 VSS.n5123 VSS.n498 585
R316 VSS.n5123 VSS.n454 585
R317 VSS.n5123 VSS.n5122 585
R318 VSS.n710 VSS.n681 585
R319 VSS.n1890 VSS.n710 585
R320 VSS.n5121 VSS.n498 585
R321 VSS.n5122 VSS.n5121 585
R322 VSS.n5121 VSS.n5120 585
R323 VSS.n686 VSS.n674 585
R324 VSS.n710 VSS.n675 585
R325 VSS.n671 VSS.n670 585
R326 VSS.n4555 VSS.n671 585
R327 VSS.n4781 VSS.n671 585
R328 VSS.n4682 VSS.n674 585
R329 VSS.n710 VSS.n673 585
R330 VSS.n4780 VSS.n670 585
R331 VSS.n4781 VSS.n4780 585
R332 VSS.n4780 VSS.n4779 585
R333 VSS.n4779 VSS.n596 585
R334 VSS.n5065 VSS.n5064 585
R335 VSS.n5065 VSS.n585 585
R336 VSS.n5063 VSS.n586 585
R337 VSS.n5059 VSS.n586 585
R338 VSS.n5062 VSS.n5061 585
R339 VSS.n5061 VSS.n5060 585
R340 VSS.n588 VSS.n587 585
R341 VSS.n5058 VSS.n588 585
R342 VSS.n5056 VSS.n5055 585
R343 VSS.n5057 VSS.n5056 585
R344 VSS.n5054 VSS.n589 585
R345 VSS.n5050 VSS.n589 585
R346 VSS.n5053 VSS.n5052 585
R347 VSS.n5052 VSS.n5051 585
R348 VSS.n591 VSS.n590 585
R349 VSS.n5049 VSS.n591 585
R350 VSS.n5047 VSS.n5046 585
R351 VSS.n5048 VSS.n5047 585
R352 VSS.n5045 VSS.n593 585
R353 VSS.n593 VSS.n592 585
R354 VSS.n5044 VSS.n5043 585
R355 VSS.n5043 VSS.n5042 585
R356 VSS.n5040 VSS.n597 585
R357 VSS.n5040 VSS.n5039 585
R358 VSS.n5034 VSS.n595 585
R359 VSS.n5038 VSS.n595 585
R360 VSS.n5036 VSS.n5035 585
R361 VSS.n5037 VSS.n5036 585
R362 VSS.n5033 VSS.n599 585
R363 VSS.n599 VSS.n598 585
R364 VSS.n5032 VSS.n5031 585
R365 VSS.n5031 VSS.n5030 585
R366 VSS.n601 VSS.n600 585
R367 VSS.n5029 VSS.n601 585
R368 VSS.n5027 VSS.n5026 585
R369 VSS.n5028 VSS.n5027 585
R370 VSS.n5025 VSS.n602 585
R371 VSS.n5021 VSS.n602 585
R372 VSS.n5024 VSS.n5023 585
R373 VSS.n5023 VSS.n5022 585
R374 VSS.n604 VSS.n603 585
R375 VSS.n5020 VSS.n604 585
R376 VSS.n5018 VSS.n5017 585
R377 VSS.n5019 VSS.n5018 585
R378 VSS.n3894 VSS.n3893 585
R379 VSS.n3895 VSS.n244 585
R380 VSS.n3894 VSS.n898 585
R381 VSS.n3894 VSS.n896 585
R382 VSS.n3895 VSS.n898 585
R383 VSS.n4503 VSS.n4502 585
R384 VSS.n4502 VSS.n4501 585
R385 VSS.n4444 VSS.n4439 585
R386 VSS.n4439 VSS.n4438 585
R387 VSS.n4510 VSS.n4509 585
R388 VSS.n4511 VSS.n4510 585
R389 VSS.n4440 VSS.n4436 585
R390 VSS.n4512 VSS.n4436 585
R391 VSS.n4515 VSS.n4514 585
R392 VSS.n4514 VSS.n4513 585
R393 VSS.n4435 VSS.n4433 585
R394 VSS.n4437 VSS.n4435 585
R395 VSS.n4520 VSS.n4430 585
R396 VSS.n4430 VSS.n4429 585
R397 VSS.n4525 VSS.n4524 585
R398 VSS.n4526 VSS.n4525 585
R399 VSS.n4431 VSS.n895 585
R400 VSS.n4527 VSS.n895 585
R401 VSS.n4530 VSS.n4529 585
R402 VSS.n4529 VSS.n4528 585
R403 VSS.n894 VSS.n892 585
R404 VSS.n4428 VSS.n894 585
R405 VSS.n4426 VSS.n4425 585
R406 VSS.n4427 VSS.n4426 585
R407 VSS.n4500 VSS.n4499 585
R408 VSS.n4497 VSS.n406 585
R409 VSS.n4499 VSS.n785 585
R410 VSS.n4499 VSS.n783 585
R411 VSS.n4497 VSS.n785 585
R412 VSS.n4650 VSS.n737 585
R413 VSS.n4650 VSS.n4649 585
R414 VSS.n741 VSS.n735 585
R415 VSS.n4647 VSS.n735 585
R416 VSS.n4645 VSS.n4644 585
R417 VSS.n4646 VSS.n4645 585
R418 VSS.n4613 VSS.n739 585
R419 VSS.n739 VSS.n738 585
R420 VSS.n4621 VSS.n4620 585
R421 VSS.n4620 VSS.n4619 585
R422 VSS.n4617 VSS.n4612 585
R423 VSS.n4618 VSS.n4617 585
R424 VSS.n4626 VSS.n4609 585
R425 VSS.n4609 VSS.n4608 585
R426 VSS.n4631 VSS.n4630 585
R427 VSS.n4632 VSS.n4631 585
R428 VSS.n4610 VSS.n782 585
R429 VSS.n4633 VSS.n782 585
R430 VSS.n4636 VSS.n4635 585
R431 VSS.n4635 VSS.n4634 585
R432 VSS.n781 VSS.n779 585
R433 VSS.n4607 VSS.n781 585
R434 VSS.n4605 VSS.n4604 585
R435 VSS.n4606 VSS.n4605 585
R436 VSS.n4648 VSS.n720 585
R437 VSS.n4657 VSS.n674 585
R438 VSS.n4656 VSS.n720 585
R439 VSS.n4652 VSS.n720 585
R440 VSS.n4657 VSS.n4656 585
R441 VSS.n5072 VSS.n5071 585
R442 VSS.n5071 VSS.n5070 585
R443 VSS.n581 VSS.n576 585
R444 VSS.n576 VSS.n575 585
R445 VSS.n5079 VSS.n5078 585
R446 VSS.n5080 VSS.n5079 585
R447 VSS.n577 VSS.n573 585
R448 VSS.n5081 VSS.n573 585
R449 VSS.n5084 VSS.n5083 585
R450 VSS.n5083 VSS.n5082 585
R451 VSS.n572 VSS.n570 585
R452 VSS.n574 VSS.n572 585
R453 VSS.n5089 VSS.n567 585
R454 VSS.n567 VSS.n566 585
R455 VSS.n5094 VSS.n5093 585
R456 VSS.n5095 VSS.n5094 585
R457 VSS.n568 VSS.n564 585
R458 VSS.n5096 VSS.n564 585
R459 VSS.n5099 VSS.n5098 585
R460 VSS.n5098 VSS.n5097 585
R461 VSS.n563 VSS.n561 585
R462 VSS.n565 VSS.n563 585
R463 VSS.n4655 VSS.n4654 585
R464 VSS.n4654 VSS.n4653 585
R465 VSS.n5069 VSS.n584 585
R466 VSS.n5068 VSS.n5067 585
R467 VSS.n3996 VSS.n3995 585
R468 VSS.n1215 VSS.n1214 585
R469 VSS.n1213 VSS.n1203 585
R470 VSS.n1207 VSS.n1204 585
R471 VSS.n1209 VSS.n1208 585
R472 VSS.n1206 VSS.n1205 585
R473 VSS.n1268 VSS.n1242 585
R474 VSS.n3962 VSS.n1242 585
R475 VSS.n3965 VSS.n3964 585
R476 VSS.n3964 VSS.n3963 585
R477 VSS.n1237 VSS.n1233 585
R478 VSS.n1233 VSS.n1232 585
R479 VSS.n3972 VSS.n3971 585
R480 VSS.n3973 VSS.n3972 585
R481 VSS.n1235 VSS.n1231 585
R482 VSS.n3974 VSS.n1231 585
R483 VSS.n3977 VSS.n3976 585
R484 VSS.n3976 VSS.n3975 585
R485 VSS.n1230 VSS.n1228 585
R486 VSS.n1230 VSS.n1229 585
R487 VSS.n1224 VSS.n1221 585
R488 VSS.n1221 VSS.n1220 585
R489 VSS.n3985 VSS.n3984 585
R490 VSS.n3986 VSS.n3985 585
R491 VSS.n1222 VSS.n1218 585
R492 VSS.n3987 VSS.n1218 585
R493 VSS.n3990 VSS.n3989 585
R494 VSS.n3989 VSS.n3988 585
R495 VSS.n3992 VSS.n1201 585
R496 VSS.n1201 VSS.n1200 585
R497 VSS.n3924 VSS.n1294 585
R498 VSS.n1294 VSS.n1293 585
R499 VSS.n3927 VSS.n3926 585
R500 VSS.n3928 VSS.n3927 585
R501 VSS.n1295 VSS.n1290 585
R502 VSS.n3929 VSS.n1290 585
R503 VSS.n3932 VSS.n3931 585
R504 VSS.n3931 VSS.n3930 585
R505 VSS.n1289 VSS.n1287 585
R506 VSS.n1292 VSS.n1289 585
R507 VSS.n1283 VSS.n1282 585
R508 VSS.n1291 VSS.n1282 585
R509 VSS.n3940 VSS.n3939 585
R510 VSS.n3944 VSS.n3940 585
R511 VSS.n3947 VSS.n3946 585
R512 VSS.n3946 VSS.n3945 585
R513 VSS.n1281 VSS.n1279 585
R514 VSS.n3943 VSS.n1281 585
R515 VSS.n3941 VSS.n1275 585
R516 VSS.n3942 VSS.n3941 585
R517 VSS.n3954 VSS.n1273 585
R518 VSS.n1273 VSS.n1272 585
R519 VSS.n3957 VSS.n3956 585
R520 VSS.n3958 VSS.n3957 585
R521 VSS.n3961 VSS.n3960 585
R522 VSS.n3960 VSS.n1271 585
R523 VSS.n3960 VSS.n3959 585
R524 VSS.n4019 VSS.n4018 585
R525 VSS.n4020 VSS.n4019 585
R526 VSS.n4019 VSS.n1126 585
R527 VSS.n3757 VSS.n3711 585
R528 VSS.n3757 VSS.n3710 585
R529 VSS.n3757 VSS.n3756 585
R530 VSS.n3710 VSS.n3709 585
R531 VSS.n3588 VSS.n3582 585
R532 VSS.n960 VSS.n958 585
R533 VSS.n4403 VSS.n960 585
R534 VSS.n3582 VSS.n960 585
R535 VSS.n3263 VSS.n1123 585
R536 VSS.n4020 VSS.n1123 585
R537 VSS.n3833 VSS.n1123 585
R538 VSS.n5473 VSS.n77 585
R539 VSS.n5474 VSS.n5473 585
R540 VSS.n5373 VSS.n244 585
R541 VSS.n244 VSS.n243 585
R542 VSS.n259 VSS.n244 585
R543 VSS.n250 VSS.n246 585
R544 VSS.n5372 VSS.n250 585
R545 VSS.n5373 VSS.n246 585
R546 VSS.n5373 VSS.n5372 585
R547 VSS.n246 VSS.n243 585
R548 VSS.n5372 VSS.n243 585
R549 VSS.n259 VSS.n246 585
R550 VSS.n418 VSS.n406 585
R551 VSS.n5193 VSS.n406 585
R552 VSS.n417 VSS.n406 585
R553 VSS.n5195 VSS.n406 585
R554 VSS.n5196 VSS.n418 585
R555 VSS.n5196 VSS.n5193 585
R556 VSS.n5193 VSS.n407 585
R557 VSS.n5196 VSS.n417 585
R558 VSS.n417 VSS.n407 585
R559 VSS.n5196 VSS.n5195 585
R560 VSS.n5189 VSS.n422 585
R561 VSS.n5190 VSS.n5189 585
R562 VSS.n1919 VSS.n674 585
R563 VSS.n1882 VSS.n674 585
R564 VSS.n1951 VSS.n674 585
R565 VSS.n1952 VSS.n1915 585
R566 VSS.n1915 VSS.n710 585
R567 VSS.n1952 VSS.n1919 585
R568 VSS.n1919 VSS.n710 585
R569 VSS.n1952 VSS.n1882 585
R570 VSS.n1882 VSS.n710 585
R571 VSS.n1952 VSS.n1951 585
R572 VSS.n4950 VSS.n620 585
R573 VSS.n1917 VSS.n620 585
R574 VSS.n4993 VSS.n4992 585
R575 VSS.n627 VSS.n626 585
R576 VSS.n4990 VSS.n4951 585
R577 VSS.n4987 VSS.n4951 585
R578 VSS.n4990 VSS.n4989 585
R579 VSS.n4989 VSS.n4988 585
R580 VSS.n150 VSS.n149 585
R581 VSS.n4145 VSS.n150 585
R582 VSS.n5427 VSS.n150 585
R583 VSS.n4276 VSS.n4255 585
R584 VSS.n4276 VSS.n32 585
R585 VSS.n5371 VSS.n244 585
R586 VSS.n248 VSS.n244 585
R587 VSS.n5369 VSS.n244 585
R588 VSS.n5370 VSS.n249 585
R589 VSS.n5372 VSS.n249 585
R590 VSS.n5371 VSS.n5370 585
R591 VSS.n5372 VSS.n5371 585
R592 VSS.n5370 VSS.n248 585
R593 VSS.n5372 VSS.n248 585
R594 VSS.n5370 VSS.n5369 585
R595 VSS.n1650 VSS.n406 585
R596 VSS.n1614 VSS.n406 585
R597 VSS.n1679 VSS.n406 585
R598 VSS.n1680 VSS.n1648 585
R599 VSS.n1648 VSS.n407 585
R600 VSS.n1680 VSS.n1650 585
R601 VSS.n1650 VSS.n407 585
R602 VSS.n1680 VSS.n1614 585
R603 VSS.n1614 VSS.n407 585
R604 VSS.n1680 VSS.n1679 585
R605 VSS.n2468 VSS.n1584 585
R606 VSS.n1682 VSS.n1584 585
R607 VSS.n1999 VSS.n674 585
R608 VSS.n1998 VSS.n674 585
R609 VSS.n2162 VSS.n674 585
R610 VSS.n2166 VSS.n2001 585
R611 VSS.n2166 VSS.n710 585
R612 VSS.n2001 VSS.n1999 585
R613 VSS.n1999 VSS.n710 585
R614 VSS.n2001 VSS.n1998 585
R615 VSS.n1998 VSS.n710 585
R616 VSS.n2162 VSS.n2001 585
R617 VSS.n373 VSS.n362 585
R618 VSS.n2466 VSS.n373 585
R619 VSS.n5254 VSS.n5253 585
R620 VSS.n367 VSS.n365 585
R621 VSS.n5257 VSS.n5256 585
R622 VSS.n5258 VSS.n5257 585
R623 VSS.n5256 VSS.n361 585
R624 VSS.n5259 VSS.n361 585
R625 VSS.n5365 VSS.n5364 585
R626 VSS.n5364 VSS.n5363 585
R627 VSS.n2621 VSS.n154 585
R628 VSS.n2925 VSS.n154 585
R629 VSS.n5425 VSS.n154 585
R630 VSS.n5426 VSS.n149 585
R631 VSS.n5427 VSS.n5426 585
R632 VSS.n5426 VSS.n5425 585
R633 VSS.n5375 VSS.n198 585
R634 VSS.n3347 VSS.n198 585
R635 VSS.n3836 VSS.n1345 585
R636 VSS.n3836 VSS.n3256 585
R637 VSS.n3836 VSS.n3835 585
R638 VSS.n3834 VSS.n3263 585
R639 VSS.n3834 VSS.n3833 585
R640 VSS.n3835 VSS.n3834 585
R641 VSS.n4406 VSS.n900 585
R642 VSS.n4407 VSS.n4406 585
R643 VSS.n4406 VSS.n4405 585
R644 VSS.n4404 VSS.n958 585
R645 VSS.n4404 VSS.n4403 585
R646 VSS.n4405 VSS.n4404 585
R647 VSS.n3831 VSS.n1008 585
R648 VSS.n3281 VSS.n1008 585
R649 VSS.n3334 VSS.n1008 585
R650 VSS.n1008 VSS.n983 585
R651 VSS.n1008 VSS.n1004 585
R652 VSS.n3339 VSS.n1008 585
R653 VSS.n1008 VSS.n1007 585
R654 VSS.n4225 VSS.n1008 585
R655 VSS.n4203 VSS.n1008 585
R656 VSS.n1008 VSS.n970 585
R657 VSS.n1008 VSS.n1005 585
R658 VSS.n4201 VSS.n1008 585
R659 VSS.n4399 VSS.n1008 585
R660 VSS.n1271 VSS.n1002 585
R661 VSS.n4400 VSS.n1002 585
R662 VSS.n4401 VSS.n4400 585
R663 VSS.n4400 VSS.n1003 585
R664 VSS.n3340 VSS.n3334 585
R665 VSS.n3340 VSS.n983 585
R666 VSS.n4400 VSS.n983 585
R667 VSS.n3340 VSS.n1004 585
R668 VSS.n4400 VSS.n1004 585
R669 VSS.n3340 VSS.n3339 585
R670 VSS.n4203 VSS.n304 585
R671 VSS.n970 VSS.n304 585
R672 VSS.n4400 VSS.n970 585
R673 VSS.n1005 VSS.n304 585
R674 VSS.n4400 VSS.n1005 585
R675 VSS.n4201 VSS.n304 585
R676 VSS.n4398 VSS.n964 585
R677 VSS.n4400 VSS.n964 585
R678 VSS.n4399 VSS.n4398 585
R679 VSS.n4400 VSS.n4399 585
R680 VSS.n4065 VSS.n6 585
R681 VSS.n6 VSS.n4 585
R682 VSS.n4069 VSS.n4067 585
R683 VSS.n4071 VSS.n4069 585
R684 VSS.n4101 VSS.n4100 585
R685 VSS.n4100 VSS.n4099 585
R686 VSS.n4074 VSS.n4070 585
R687 VSS.n4098 VSS.n4070 585
R688 VSS.n4096 VSS.n4095 585
R689 VSS.n4097 VSS.n4096 585
R690 VSS.n4078 VSS.n4073 585
R691 VSS.n4073 VSS.n4072 585
R692 VSS.n4090 VSS.n4089 585
R693 VSS.n4089 VSS.n4088 585
R694 VSS.n4085 VSS.n4084 585
R695 VSS.n4087 VSS.n4085 585
R696 VSS.n4080 VSS.n1015 585
R697 VSS.n4086 VSS.n1015 585
R698 VSS.n4324 VSS.n4323 585
R699 VSS.n4325 VSS.n4324 585
R700 VSS.n1017 VSS.n1014 585
R701 VSS.n4326 VSS.n1014 585
R702 VSS.n4329 VSS.n4328 585
R703 VSS.n4328 VSS.n4327 585
R704 VSS.n4397 VSS.n4396 585
R705 VSS.n4396 VSS.n4395 585
R706 VSS.n4336 VSS.n4333 585
R707 VSS.n4394 VSS.n4333 585
R708 VSS.n4392 VSS.n4391 585
R709 VSS.n4393 VSS.n4392 585
R710 VSS.n4338 VSS.n4335 585
R711 VSS.n4335 VSS.n4334 585
R712 VSS.n4364 VSS.n4363 585
R713 VSS.n4363 VSS.n4362 585
R714 VSS.n4360 VSS.n4359 585
R715 VSS.n4361 VSS.n4360 585
R716 VSS.n4342 VSS.n4341 585
R717 VSS.n4350 VSS.n4341 585
R718 VSS.n4353 VSS.n4352 585
R719 VSS.n4352 VSS.n4351 585
R720 VSS.n4349 VSS.n4348 585
R721 VSS.n4349 VSS.n338 585
R722 VSS.n336 VSS.n334 585
R723 VSS.n5289 VSS.n336 585
R724 VSS.n5293 VSS.n5292 585
R725 VSS.n5292 VSS.n5291 585
R726 VSS.n1517 VSS.n337 585
R727 VSS.n5290 VSS.n337 585
R728 VSS.n1523 VSS.n1522 585
R729 VSS.n1524 VSS.n1523 585
R730 VSS.n1491 VSS.n1489 585
R731 VSS.n1525 VSS.n1491 585
R732 VSS.n2560 VSS.n2559 585
R733 VSS.n2559 VSS.n2558 585
R734 VSS.n1528 VSS.n1492 585
R735 VSS.n2557 VSS.n1492 585
R736 VSS.n2555 VSS.n2554 585
R737 VSS.n2556 VSS.n2555 585
R738 VSS.n1532 VSS.n1527 585
R739 VSS.n1527 VSS.n1526 585
R740 VSS.n2549 VSS.n2548 585
R741 VSS.n2548 VSS.n2547 585
R742 VSS.n1537 VSS.n1534 585
R743 VSS.n2546 VSS.n1534 585
R744 VSS.n2544 VSS.n2543 585
R745 VSS.n2545 VSS.n2544 585
R746 VSS.n1541 VSS.n1536 585
R747 VSS.n1536 VSS.n1535 585
R748 VSS.n2538 VSS.n2537 585
R749 VSS.n2537 VSS.n2536 585
R750 VSS.n2535 VSS.n2534 585
R751 VSS.n2535 VSS.n342 585
R752 VSS.n2529 VSS.n2528 585
R753 VSS.n2528 VSS.n2527 585
R754 VSS.n1566 VSS.n1563 585
R755 VSS.n2526 VSS.n1563 585
R756 VSS.n2524 VSS.n2523 585
R757 VSS.n2525 VSS.n2524 585
R758 VSS.n1568 VSS.n1565 585
R759 VSS.n1565 VSS.n1564 585
R760 VSS.n2236 VSS.n2235 585
R761 VSS.n2235 VSS.n2234 585
R762 VSS.n2231 VSS.n2230 585
R763 VSS.n2233 VSS.n2230 585
R764 VSS.n2244 VSS.n2243 585
R765 VSS.n2245 VSS.n2244 585
R766 VSS.n2248 VSS.n2247 585
R767 VSS.n2247 VSS.n2246 585
R768 VSS.n2249 VSS.n2225 585
R769 VSS.n2225 VSS.n2224 585
R770 VSS.n2285 VSS.n2284 585
R771 VSS.n2286 VSS.n2285 585
R772 VSS.n2227 VSS.n2223 585
R773 VSS.n2287 VSS.n2223 585
R774 VSS.n2290 VSS.n2289 585
R775 VSS.n2289 VSS.n2288 585
R776 VSS.n2296 VSS.n2295 585
R777 VSS.n2296 VSS.n346 585
R778 VSS.n2299 VSS.n2298 585
R779 VSS.n2298 VSS.n2297 585
R780 VSS.n2300 VSS.n2127 585
R781 VSS.n2127 VSS.n2126 585
R782 VSS.n2309 VSS.n2308 585
R783 VSS.n2310 VSS.n2309 585
R784 VSS.n2130 VSS.n2125 585
R785 VSS.n2311 VSS.n2125 585
R786 VSS.n2313 VSS.n2124 585
R787 VSS.n2313 VSS.n2312 585
R788 VSS.n2316 VSS.n2315 585
R789 VSS.n2315 VSS.n2314 585
R790 VSS.n2121 VSS.n2120 585
R791 VSS.n2120 VSS.n2119 585
R792 VSS.n2326 VSS.n2325 585
R793 VSS.n2327 VSS.n2326 585
R794 VSS.n2118 VSS.n2115 585
R795 VSS.n2328 VSS.n2118 585
R796 VSS.n2331 VSS.n2330 585
R797 VSS.n2330 VSS.n2329 585
R798 VSS.n2116 VSS.n349 585
R799 VSS.n349 VSS.n347 585
R800 VSS.n1198 VSS.n1197 585
R801 VSS.n3998 VSS.n1198 585
R802 VSS.n4001 VSS.n4000 585
R803 VSS.n4000 VSS.n3999 585
R804 VSS.n4002 VSS.n1195 585
R805 VSS.n1195 VSS.n1193 585
R806 VSS.n4004 VSS.n4003 585
R807 VSS.n4005 VSS.n4004 585
R808 VSS.n1196 VSS.n1194 585
R809 VSS.n1194 VSS.n1192 585
R810 VSS.n3755 VSS.n3754 585
R811 VSS.n3754 VSS.n3753 585
R812 VSS.n3750 VSS.n3749 585
R813 VSS.n3751 VSS.n3750 585
R814 VSS.n3748 VSS.n3747 585
R815 VSS.n3747 VSS.n3712 585
R816 VSS.n3746 VSS.n3713 585
R817 VSS.n3746 VSS.n3745 585
R818 VSS.n3740 VSS.n3714 585
R819 VSS.n3744 VSS.n3714 585
R820 VSS.n3742 VSS.n3741 585
R821 VSS.n3743 VSS.n3742 585
R822 VSS.n3739 VSS.n3715 585
R823 VSS.n3735 VSS.n3715 585
R824 VSS.n3738 VSS.n3737 585
R825 VSS.n3737 VSS.n3736 585
R826 VSS.n3717 VSS.n3716 585
R827 VSS.n3734 VSS.n3717 585
R828 VSS.n3732 VSS.n3731 585
R829 VSS.n3733 VSS.n3732 585
R830 VSS.n3730 VSS.n3719 585
R831 VSS.n3719 VSS.n3718 585
R832 VSS.n3729 VSS.n3728 585
R833 VSS.n3728 VSS.n3727 585
R834 VSS.n3721 VSS.n3720 585
R835 VSS.n3726 VSS.n3721 585
R836 VSS.n3724 VSS.n3723 585
R837 VSS.n3725 VSS.n3724 585
R838 VSS.n4017 VSS.n4016 585
R839 VSS.n4016 VSS.n4015 585
R840 VSS.n1146 VSS.n1127 585
R841 VSS.n1146 VSS.n1128 585
R842 VSS.n1149 VSS.n1148 585
R843 VSS.n1148 VSS.n1147 585
R844 VSS.n1151 VSS.n1150 585
R845 VSS.n1152 VSS.n1151 585
R846 VSS.n1144 VSS.n1143 585
R847 VSS.n1153 VSS.n1144 585
R848 VSS.n1156 VSS.n1155 585
R849 VSS.n1155 VSS.n1154 585
R850 VSS.n1157 VSS.n1131 585
R851 VSS.n1145 VSS.n1131 585
R852 VSS.n1159 VSS.n1158 585
R853 VSS.n1160 VSS.n1159 585
R854 VSS.n1142 VSS.n1130 585
R855 VSS.n1130 VSS.n1129 585
R856 VSS.n1141 VSS.n1140 585
R857 VSS.n1140 VSS.n1139 585
R858 VSS.n1133 VSS.n1132 585
R859 VSS.n1138 VSS.n1133 585
R860 VSS.n1137 VSS.n1136 585
R861 VSS.n1134 VSS.n74 585
R862 VSS.n5476 VSS.n71 585
R863 VSS.n5477 VSS.n5476 585
R864 VSS.n72 VSS.n71 585
R865 VSS.n5478 VSS.n72 585
R866 VSS.n5481 VSS.n5480 585
R867 VSS.n5480 VSS.n5479 585
R868 VSS.n5482 VSS.n70 585
R869 VSS.n70 VSS.n69 585
R870 VSS.n5484 VSS.n5483 585
R871 VSS.n5485 VSS.n5484 585
R872 VSS.n67 VSS.n66 585
R873 VSS.n5486 VSS.n67 585
R874 VSS.n5489 VSS.n5488 585
R875 VSS.n5488 VSS.n5487 585
R876 VSS.n5490 VSS.n65 585
R877 VSS.n68 VSS.n65 585
R878 VSS.n5492 VSS.n5491 585
R879 VSS.n5493 VSS.n5492 585
R880 VSS.n63 VSS.n62 585
R881 VSS.n5494 VSS.n63 585
R882 VSS.n5497 VSS.n5496 585
R883 VSS.n5496 VSS.n5495 585
R884 VSS.n5498 VSS.n60 585
R885 VSS.n64 VSS.n60 585
R886 VSS.n5500 VSS.n5499 585
R887 VSS.n5501 VSS.n5500 585
R888 VSS.n5514 VSS.n5513 585
R889 VSS.n5513 VSS.n5512 585
R890 VSS.n5515 VSS.n44 585
R891 VSS.n44 VSS.n43 585
R892 VSS.n5517 VSS.n5516 585
R893 VSS.n5518 VSS.n5517 585
R894 VSS.n42 VSS.n41 585
R895 VSS.n5519 VSS.n42 585
R896 VSS.n5522 VSS.n5521 585
R897 VSS.n5521 VSS.n5520 585
R898 VSS.n5523 VSS.n40 585
R899 VSS.n40 VSS.n39 585
R900 VSS.n5525 VSS.n5524 585
R901 VSS.n5526 VSS.n5525 585
R902 VSS.n37 VSS.n36 585
R903 VSS.n5527 VSS.n37 585
R904 VSS.n5530 VSS.n5529 585
R905 VSS.n5529 VSS.n5528 585
R906 VSS.n5531 VSS.n35 585
R907 VSS.n38 VSS.n35 585
R908 VSS.n5533 VSS.n5532 585
R909 VSS.n5533 VSS.n34 585
R910 VSS.n5535 VSS.n5534 585
R911 VSS.n5537 VSS.n5536 585
R912 VSS.n5539 VSS.n28 585
R913 VSS.n5540 VSS.n5539 585
R914 VSS.n29 VSS.n28 585
R915 VSS.n5541 VSS.n29 585
R916 VSS.n5544 VSS.n5543 585
R917 VSS.n5543 VSS.n5542 585
R918 VSS.n5545 VSS.n27 585
R919 VSS.n30 VSS.n27 585
R920 VSS.n5547 VSS.n5546 585
R921 VSS.n5548 VSS.n5547 585
R922 VSS.n13 VSS.n12 585
R923 VSS.n5549 VSS.n13 585
R924 VSS.n5552 VSS.n5551 585
R925 VSS.n5551 VSS.n5550 585
R926 VSS.n5553 VSS.n10 585
R927 VSS.n14 VSS.n10 585
R928 VSS.n5555 VSS.n5554 585
R929 VSS.n5556 VSS.n5555 585
R930 VSS.n11 VSS.n8 585
R931 VSS.n5557 VSS.n8 585
R932 VSS.n5559 VSS.n9 585
R933 VSS.n5559 VSS.n5558 585
R934 VSS.n5560 VSS.n5 585
R935 VSS.n5563 VSS.n5562 585
R936 VSS.n1185 VSS.n1184 584.309
R937 VSS.n5283 VSS.n5282 568.683
R938 VSS.n1211 VSS.n1199 558.078
R939 VSS.n4012 VSS.n1163 522.542
R940 VSS.t104 VSS.t0 519.213
R941 VSS.t0 VSS.t48 519.213
R942 VSS.t48 VSS.t30 519.213
R943 VSS.t30 VSS.t40 519.213
R944 VSS.t40 VSS.t18 519.213
R945 VSS.t28 VSS.t22 519.213
R946 VSS.t22 VSS.t35 519.213
R947 VSS.t35 VSS.t1 519.213
R948 VSS.t1 VSS.t36 519.213
R949 VSS.n4011 VSS.n1165 493.93
R950 VSS.n5289 VSS.n5288 466.325
R951 VSS.n5016 VSS.n607 426.668
R952 VSS.n4088 VSS.t54 353.505
R953 VSS.n4350 VSS.t60 353.505
R954 VSS.n2547 VSS.t69 353.505
R955 VSS.n2245 VSS.t57 353.505
R956 VSS.n2314 VSS.t72 353.505
R957 VSS.n4548 VSS.t69 346.457
R958 VSS.n3053 VSS.t69 346.457
R959 VSS.n3115 VSS.t69 346.457
R960 VSS.n3082 VSS.t69 346.457
R961 VSS.n340 VSS.t28 346.142
R962 VSS.n4276 VSS.t54 331.916
R963 VSS.n5473 VSS.t54 331.916
R964 VSS.n3582 VSS.t54 331.916
R965 VSS.n3796 VSS.t54 331.916
R966 VSS.n1063 VSS.t54 331.916
R967 VSS.t72 VSS.n373 128.062
R968 VSS.n5229 VSS.t72 128.062
R969 VSS.t72 VSS.n620 128.062
R970 VSS.n5120 VSS.t72 128.062
R971 VSS.n4779 VSS.t72 128.062
R972 VSS.n4072 VSS.t54 323.42
R973 VSS.n4361 VSS.t60 323.42
R974 VSS.n1526 VSS.t69 323.42
R975 VSS.n2233 VSS.t57 323.42
R976 VSS.n2312 VSS.t72 323.42
R977 VSS.n4307 VSS.t54 319.149
R978 VSS.n5455 VSS.t54 319.149
R979 VSS.n3710 VSS.t54 319.149
R980 VSS.n4020 VSS.t54 319.149
R981 VSS.n4145 VSS.t54 319.149
R982 VSS.n2357 VSS.t72 130.675
R983 VSS.t72 VSS.n374 130.675
R984 VSS.n4948 VSS.t72 130.675
R985 VSS.t72 VSS.n621 130.675
R986 VSS.n4740 VSS.t72 130.675
R987 VSS.n367 VSS.t72 302.586
R988 VSS.n4964 VSS.t72 302.586
R989 VSS.n626 VSS.t72 302.586
R990 VSS.n613 VSS.t72 302.586
R991 VSS.n5042 VSS.t72 302.586
R992 VSS.n5284 VSS.n346 300.856
R993 VSS.n4660 VSS.n4659 292.5
R994 VSS.n1895 VSS.n1888 292.5
R995 VSS.n1949 VSS.n1880 292.5
R996 VSS.n2180 VSS.n2179 292.5
R997 VSS.n4662 VSS.n4661 292.5
R998 VSS.n4664 VSS.n716 292.5
R999 VSS.n4666 VSS.n715 292.5
R1000 VSS.n4669 VSS.n4668 292.5
R1001 VSS.n4671 VSS.n4670 292.5
R1002 VSS.n4673 VSS.n713 292.5
R1003 VSS.n4675 VSS.n712 292.5
R1004 VSS.n4678 VSS.n4677 292.5
R1005 VSS.n1897 VSS.n1887 292.5
R1006 VSS.n1900 VSS.n1899 292.5
R1007 VSS.n1902 VSS.n1901 292.5
R1008 VSS.n1904 VSS.n1885 292.5
R1009 VSS.n1906 VSS.n1884 292.5
R1010 VSS.n1909 VSS.n1908 292.5
R1011 VSS.n1911 VSS.n1910 292.5
R1012 VSS.n1913 VSS.n1881 292.5
R1013 VSS.n1947 VSS.n1946 292.5
R1014 VSS.n1945 VSS.n1944 292.5
R1015 VSS.n1942 VSS.n1921 292.5
R1016 VSS.n1940 VSS.n1939 292.5
R1017 VSS.n1938 VSS.n1937 292.5
R1018 VSS.n1935 VSS.n1923 292.5
R1019 VSS.n1933 VSS.n1932 292.5
R1020 VSS.n1931 VSS.n1930 292.5
R1021 VSS.n2182 VSS.n2181 292.5
R1022 VSS.n2184 VSS.n2171 292.5
R1023 VSS.n2186 VSS.n2170 292.5
R1024 VSS.n2189 VSS.n2188 292.5
R1025 VSS.n2191 VSS.n2190 292.5
R1026 VSS.n2193 VSS.n2168 292.5
R1027 VSS.n2195 VSS.n2164 292.5
R1028 VSS.n2198 VSS.n2197 292.5
R1029 VSS.n2201 VSS.n2200 292.5
R1030 VSS.n2203 VSS.n2160 292.5
R1031 VSS.n2206 VSS.n2205 292.5
R1032 VSS.n2208 VSS.n2207 292.5
R1033 VSS.n2210 VSS.n2158 292.5
R1034 VSS.n2212 VSS.n2157 292.5
R1035 VSS.n2215 VSS.n2214 292.5
R1036 VSS.n2217 VSS.n2216 292.5
R1037 VSS.n2219 VSS.n2155 292.5
R1038 VSS.n3085 VSS.n3084 292.5
R1039 VSS.n3084 VSS.n3083 292.5
R1040 VSS.n1448 VSS.n1444 292.5
R1041 VSS.n3081 VSS.n1444 292.5
R1042 VSS.n3079 VSS.n3078 292.5
R1043 VSS.n3080 VSS.n3079 292.5
R1044 VSS.n2943 VSS.n1446 292.5
R1045 VSS.n1446 VSS.n1445 292.5
R1046 VSS.n2941 VSS.n2931 292.5
R1047 VSS.n2931 VSS.n2930 292.5
R1048 VSS.n2958 VSS.n2957 292.5
R1049 VSS.n2959 VSS.n2958 292.5
R1050 VSS.n2937 VSS.n2592 292.5
R1051 VSS.n2960 VSS.n2592 292.5
R1052 VSS.n2963 VSS.n2962 292.5
R1053 VSS.n2962 VSS.n2961 292.5
R1054 VSS.n2591 VSS.n2586 292.5
R1055 VSS.n2929 VSS.n2591 292.5
R1056 VSS.n2927 VSS.n2585 292.5
R1057 VSS.n3082 VSS.n404 292.5
R1058 VSS.n2393 VSS.n2392 292.5
R1059 VSS.n2401 VSS.n2400 292.5
R1060 VSS.n2404 VSS.n2403 292.5
R1061 VSS.n2055 VSS.n2054 292.5
R1062 VSS.n2052 VSS.n2051 292.5
R1063 VSS.n2416 VSS.n2415 292.5
R1064 VSS.n2419 VSS.n2418 292.5
R1065 VSS.n2042 VSS.n2041 292.5
R1066 VSS.n2039 VSS.n2038 292.5
R1067 VSS.n2431 VSS.n2430 292.5
R1068 VSS.n1928 VSS.n1925 292.5
R1069 VSS.n1926 VSS.n393 292.5
R1070 VSS.n2175 VSS.n2174 292.5
R1071 VSS.n2177 VSS.n2173 292.5
R1072 VSS.n1705 VSS.n1704 292.5
R1073 VSS.n1796 VSS.n1703 292.5
R1074 VSS.n1799 VSS.n1798 292.5
R1075 VSS.n1793 VSS.n1792 292.5
R1076 VSS.n1717 VSS.n1714 292.5
R1077 VSS.n1716 VSS.n1715 292.5
R1078 VSS.n1779 VSS.n1778 292.5
R1079 VSS.n1773 VSS.n1772 292.5
R1080 VSS.n1721 VSS.n1720 292.5
R1081 VSS.n1723 VSS.n1722 292.5
R1082 VSS.n3158 VSS.n3157 292.5
R1083 VSS.n3152 VSS.n3151 292.5
R1084 VSS.n1412 VSS.n1407 292.5
R1085 VSS.n3147 VSS.n3146 292.5
R1086 VSS.n2756 VSS.n1410 292.5
R1087 VSS.n2754 VSS.n2753 292.5
R1088 VSS.n2766 VSS.n2765 292.5
R1089 VSS.n2747 VSS.n2746 292.5
R1090 VSS.n2773 VSS.n2772 292.5
R1091 VSS.n2745 VSS.n2744 292.5
R1092 VSS.n4559 VSS.n4558 292.5
R1093 VSS.n836 VSS.n814 292.5
R1094 VSS.n834 VSS.n813 292.5
R1095 VSS.n4569 VSS.n4568 292.5
R1096 VSS.n4572 VSS.n4571 292.5
R1097 VSS.n803 VSS.n799 292.5
R1098 VSS.n801 VSS.n798 292.5
R1099 VSS.n4582 VSS.n4581 292.5
R1100 VSS.n4585 VSS.n4584 292.5
R1101 VSS.n4552 VSS.n4551 292.5
R1102 VSS.n4549 VSS.n4548 292.5
R1103 VSS.n4445 VSS.n841 292.5
R1104 VSS.n4547 VSS.n841 292.5
R1105 VSS.n4545 VSS.n4544 292.5
R1106 VSS.n4546 VSS.n4545 292.5
R1107 VSS.n922 VSS.n843 292.5
R1108 VSS.n843 VSS.n842 292.5
R1109 VSS.n928 VSS.n927 292.5
R1110 VSS.n929 VSS.n928 292.5
R1111 VSS.n932 VSS.n931 292.5
R1112 VSS.n931 VSS.n930 292.5
R1113 VSS.n914 VSS.n910 292.5
R1114 VSS.n914 VSS.n913 292.5
R1115 VSS.n909 VSS.n904 292.5
R1116 VSS.n912 VSS.n904 292.5
R1117 VSS.n942 VSS.n941 292.5
R1118 VSS.n942 VSS.n903 292.5
R1119 VSS.n943 VSS.n868 292.5
R1120 VSS.n944 VSS.n943 292.5
R1121 VSS.n902 VSS.n867 292.5
R1122 VSS.n3921 VSS.n3920 292.5
R1123 VSS.n3918 VSS.n3917 292.5
R1124 VSS.n3916 VSS.n3915 292.5
R1125 VSS.n3913 VSS.n3912 292.5
R1126 VSS.n3911 VSS.n3910 292.5
R1127 VSS.n3908 VSS.n3907 292.5
R1128 VSS.n3906 VSS.n3905 292.5
R1129 VSS.n3903 VSS.n3902 292.5
R1130 VSS.n3901 VSS.n3900 292.5
R1131 VSS.n3898 VSS.n3897 292.5
R1132 VSS.n949 VSS.n947 292.5
R1133 VSS.n3225 VSS.n266 292.5
R1134 VSS.n3228 VSS.n3227 292.5
R1135 VSS.n3230 VSS.n3229 292.5
R1136 VSS.n3233 VSS.n3232 292.5
R1137 VSS.n3235 VSS.n3234 292.5
R1138 VSS.n3238 VSS.n3237 292.5
R1139 VSS.n3240 VSS.n3239 292.5
R1140 VSS.n3243 VSS.n3242 292.5
R1141 VSS.n3245 VSS.n3244 292.5
R1142 VSS.n3248 VSS.n3247 292.5
R1143 VSS.n3250 VSS.n3249 292.5
R1144 VSS.n3253 VSS.n3252 292.5
R1145 VSS.n3255 VSS.n3254 292.5
R1146 VSS.n2870 VSS.n279 292.5
R1147 VSS.n2873 VSS.n2872 292.5
R1148 VSS.n2875 VSS.n2874 292.5
R1149 VSS.n2878 VSS.n2877 292.5
R1150 VSS.n2880 VSS.n2879 292.5
R1151 VSS.n2883 VSS.n2882 292.5
R1152 VSS.n2885 VSS.n2884 292.5
R1153 VSS.n2888 VSS.n2887 292.5
R1154 VSS.n2890 VSS.n2889 292.5
R1155 VSS.n2893 VSS.n2892 292.5
R1156 VSS.n2896 VSS.n2895 292.5
R1157 VSS.n2899 VSS.n2898 292.5
R1158 VSS.n2902 VSS.n2901 292.5
R1159 VSS.n2904 VSS.n2903 292.5
R1160 VSS.n2907 VSS.n2906 292.5
R1161 VSS.n2909 VSS.n2908 292.5
R1162 VSS.n2912 VSS.n2911 292.5
R1163 VSS.n2914 VSS.n2913 292.5
R1164 VSS.n2917 VSS.n2916 292.5
R1165 VSS.n2919 VSS.n2918 292.5
R1166 VSS.n2922 VSS.n2921 292.5
R1167 VSS.n2924 VSS.n2923 292.5
R1168 VSS.n2620 VSS.n285 292.5
R1169 VSS.n2619 VSS.n2618 292.5
R1170 VSS.n2616 VSS.n2615 292.5
R1171 VSS.n2613 VSS.n2612 292.5
R1172 VSS.n2611 VSS.n2610 292.5
R1173 VSS.n2608 VSS.n2607 292.5
R1174 VSS.n2606 VSS.n2605 292.5
R1175 VSS.n2603 VSS.n2602 292.5
R1176 VSS.n2601 VSS.n2600 292.5
R1177 VSS.n2598 VSS.n2597 292.5
R1178 VSS.n2596 VSS.n2595 292.5
R1179 VSS.n1495 VSS.n1494 292.5
R1180 VSS.n1498 VSS.n1497 292.5
R1181 VSS.n1500 VSS.n1499 292.5
R1182 VSS.n1503 VSS.n1502 292.5
R1183 VSS.n1505 VSS.n1504 292.5
R1184 VSS.n1508 VSS.n1507 292.5
R1185 VSS.n1510 VSS.n1509 292.5
R1186 VSS.n1513 VSS.n1512 292.5
R1187 VSS.n1516 VSS.n1515 292.5
R1188 VSS.n4495 VSS.n4494 292.5
R1189 VSS.n4492 VSS.n4491 292.5
R1190 VSS.n4489 VSS.n4465 292.5
R1191 VSS.n4487 VSS.n4486 292.5
R1192 VSS.n4485 VSS.n4484 292.5
R1193 VSS.n4482 VSS.n4467 292.5
R1194 VSS.n4480 VSS.n4479 292.5
R1195 VSS.n4478 VSS.n4477 292.5
R1196 VSS.n4475 VSS.n4469 292.5
R1197 VSS.n4473 VSS.n4472 292.5
R1198 VSS.n4470 VSS.n840 292.5
R1199 VSS.n3189 VSS.n3188 292.5
R1200 VSS.n3191 VSS.n3190 292.5
R1201 VSS.n3193 VSS.n3186 292.5
R1202 VSS.n3195 VSS.n3185 292.5
R1203 VSS.n3198 VSS.n3197 292.5
R1204 VSS.n3200 VSS.n3199 292.5
R1205 VSS.n3202 VSS.n3183 292.5
R1206 VSS.n3204 VSS.n3182 292.5
R1207 VSS.n3207 VSS.n3206 292.5
R1208 VSS.n3209 VSS.n3208 292.5
R1209 VSS.n3211 VSS.n3180 292.5
R1210 VSS.n3213 VSS.n3179 292.5
R1211 VSS.n5199 VSS.n5198 292.5
R1212 VSS.n5201 VSS.n413 292.5
R1213 VSS.n5204 VSS.n5203 292.5
R1214 VSS.n5206 VSS.n5205 292.5
R1215 VSS.n5208 VSS.n411 292.5
R1216 VSS.n5210 VSS.n410 292.5
R1217 VSS.n5213 VSS.n5212 292.5
R1218 VSS.n5215 VSS.n5214 292.5
R1219 VSS.n5217 VSS.n408 292.5
R1220 VSS.n5219 VSS.n405 292.5
R1221 VSS.n5222 VSS.n5221 292.5
R1222 VSS.n1624 VSS.n1623 292.5
R1223 VSS.n1626 VSS.n1625 292.5
R1224 VSS.n1628 VSS.n1621 292.5
R1225 VSS.n1630 VSS.n1620 292.5
R1226 VSS.n1633 VSS.n1632 292.5
R1227 VSS.n1635 VSS.n1634 292.5
R1228 VSS.n1637 VSS.n1618 292.5
R1229 VSS.n1639 VSS.n1617 292.5
R1230 VSS.n1642 VSS.n1641 292.5
R1231 VSS.n1644 VSS.n1643 292.5
R1232 VSS.n1646 VSS.n1615 292.5
R1233 VSS.n1677 VSS.n1676 292.5
R1234 VSS.n1675 VSS.n1674 292.5
R1235 VSS.n1672 VSS.n1653 292.5
R1236 VSS.n1670 VSS.n1669 292.5
R1237 VSS.n1668 VSS.n1667 292.5
R1238 VSS.n1665 VSS.n1655 292.5
R1239 VSS.n1663 VSS.n1662 292.5
R1240 VSS.n1661 VSS.n1660 292.5
R1241 VSS.n1658 VSS.n1560 292.5
R1242 VSS.n1382 VSS.n1357 292.5
R1243 VSS.n1380 VSS.n1379 292.5
R1244 VSS.n1378 VSS.n1377 292.5
R1245 VSS.n1375 VSS.n1359 292.5
R1246 VSS.n1373 VSS.n1372 292.5
R1247 VSS.n1371 VSS.n1370 292.5
R1248 VSS.n1368 VSS.n1361 292.5
R1249 VSS.n1366 VSS.n1365 292.5
R1250 VSS.n1363 VSS.n415 292.5
R1251 VSS.n3216 VSS.n3215 292.5
R1252 VSS.n1387 VSS.n1386 292.5
R1253 VSS.n1385 VSS.n1384 292.5
R1254 VSS.n5126 VSS.n5125 292.5
R1255 VSS.n496 VSS.n495 292.5
R1256 VSS.n491 VSS.n468 292.5
R1257 VSS.n489 VSS.n467 292.5
R1258 VSS.n487 VSS.n486 292.5
R1259 VSS.n5147 VSS.n5146 292.5
R1260 VSS.n5149 VSS.n455 292.5
R1261 VSS.n5152 VSS.n5151 292.5
R1262 VSS.n3217 VSS.n448 292.5
R1263 VSS.n3218 VSS.n447 292.5
R1264 VSS.n609 VSS.n503 292.5
R1265 VSS.n4880 VSS.n4879 292.5
R1266 VSS.n4872 VSS.n4871 292.5
R1267 VSS.n4869 VSS.n4868 292.5
R1268 VSS.n4863 VSS.n4862 292.5
R1269 VSS.n4860 VSS.n4859 292.5
R1270 VSS.n4850 VSS.n4849 292.5
R1271 VSS.n4847 VSS.n516 292.5
R1272 VSS.n515 VSS.n514 292.5
R1273 VSS.n5118 VSS.n5117 292.5
R1274 VSS.n4801 VSS.n508 292.5
R1275 VSS.n681 VSS.n501 292.5
R1276 VSS.n1891 VSS.n1890 292.5
R1277 VSS.n1893 VSS.n1892 292.5
R1278 VSS.n708 VSS.n707 292.5
R1279 VSS.n704 VSS.n703 292.5
R1280 VSS.n702 VSS.n701 292.5
R1281 VSS.n699 VSS.n698 292.5
R1282 VSS.n697 VSS.n696 292.5
R1283 VSS.n694 VSS.n693 292.5
R1284 VSS.n692 VSS.n691 292.5
R1285 VSS.n689 VSS.n688 292.5
R1286 VSS.n687 VSS.n686 292.5
R1287 VSS.n685 VSS.n675 292.5
R1288 VSS.n4680 VSS.n4679 292.5
R1289 VSS.n4682 VSS.n672 292.5
R1290 VSS.n705 VSS.n673 292.5
R1291 VSS.n706 VSS.n683 292.5
R1292 VSS.n4774 VSS.n596 292.5
R1293 VSS.n4777 VSS.n4776 292.5
R1294 VSS.n4769 VSS.n4690 292.5
R1295 VSS.n4732 VSS.n4724 292.5
R1296 VSS.n4735 VSS.n4725 292.5
R1297 VSS.n4734 VSS.n4727 292.5
R1298 VSS.n4738 VSS.n4726 292.5
R1299 VSS.n4737 VSS.n4728 292.5
R1300 VSS.n4743 VSS.n4742 292.5
R1301 VSS.n4731 VSS.n539 292.5
R1302 VSS.n4685 VSS.n538 292.5
R1303 VSS.n3707 VSS.n3706 292.5
R1304 VSS.n3709 VSS.n3589 292.5
R1305 VSS.n3611 VSS.n3588 292.5
R1306 VSS.n3675 VSS.n3674 292.5
R1307 VSS.n3672 VSS.n3671 292.5
R1308 VSS.n3666 VSS.n3665 292.5
R1309 VSS.n3663 VSS.n3662 292.5
R1310 VSS.n3657 VSS.n3656 292.5
R1311 VSS.n3654 VSS.n3653 292.5
R1312 VSS.n3760 VSS.n3759 292.5
R1313 VSS.n3799 VSS.n3798 292.5
R1314 VSS.n3565 VSS.n3564 292.5
R1315 VSS.n3561 VSS.n3560 292.5
R1316 VSS.n3573 VSS.n3572 292.5
R1317 VSS.n3553 VSS.n3552 292.5
R1318 VSS.n3532 VSS.n3531 292.5
R1319 VSS.n3530 VSS.n3529 292.5
R1320 VSS.n3794 VSS.n3793 292.5
R1321 VSS.n3782 VSS.n1118 292.5
R1322 VSS.n4023 VSS.n4022 292.5
R1323 VSS.n3335 VSS.n77 292.5
R1324 VSS.n5458 VSS.n5457 292.5
R1325 VSS.n5453 VSS.n5452 292.5
R1326 VSS.n118 VSS.n117 292.5
R1327 VSS.n121 VSS.n120 292.5
R1328 VSS.n128 VSS.n127 292.5
R1329 VSS.n126 VSS.n125 292.5
R1330 VSS.n114 VSS.n90 292.5
R1331 VSS.n89 VSS.n88 292.5
R1332 VSS.n5471 VSS.n5470 292.5
R1333 VSS.n4045 VSS.n82 292.5
R1334 VSS.n5474 VSS.n76 292.5
R1335 VSS.n1434 VSS.n420 292.5
R1336 VSS.n3115 VSS.n420 292.5
R1337 VSS.n1433 VSS.n1426 292.5
R1338 VSS.n3116 VSS.n1426 292.5
R1339 VSS.n3119 VSS.n3118 292.5
R1340 VSS.n3118 VSS.n3117 292.5
R1341 VSS.n1430 VSS.n1425 292.5
R1342 VSS.n3114 VSS.n1425 292.5
R1343 VSS.n3112 VSS.n3111 292.5
R1344 VSS.n3113 VSS.n3112 292.5
R1345 VSS.n2833 VSS.n1428 292.5
R1346 VSS.n1428 VSS.n1427 292.5
R1347 VSS.n2839 VSS.n2838 292.5
R1348 VSS.n2840 VSS.n2839 292.5
R1349 VSS.n2829 VSS.n2814 292.5
R1350 VSS.n2841 VSS.n2814 292.5
R1351 VSS.n2844 VSS.n2843 292.5
R1352 VSS.n2843 VSS.n2842 292.5
R1353 VSS.n2813 VSS.n2736 292.5
R1354 VSS.n2817 VSS.n2813 292.5
R1355 VSS.n2815 VSS.n2735 292.5
R1356 VSS.n2732 VSS.n242 292.5
R1357 VSS.n1955 VSS.n422 292.5
R1358 VSS.n1877 VSS.n1876 292.5
R1359 VSS.n1872 VSS.n1871 292.5
R1360 VSS.n1816 VSS.n1814 292.5
R1361 VSS.n1838 VSS.n1837 292.5
R1362 VSS.n1829 VSS.n1828 292.5
R1363 VSS.n1825 VSS.n1824 292.5
R1364 VSS.n1811 VSS.n435 292.5
R1365 VSS.n434 VSS.n433 292.5
R1366 VSS.n5187 VSS.n5186 292.5
R1367 VSS.n439 VSS.n427 292.5
R1368 VSS.n5190 VSS.n419 292.5
R1369 VSS.n4950 VSS.n628 292.5
R1370 VSS.n4831 VSS.n629 292.5
R1371 VSS.n4946 VSS.n4944 292.5
R1372 VSS.n4904 VSS.n634 292.5
R1373 VSS.n4911 VSS.n4910 292.5
R1374 VSS.n4919 VSS.n4918 292.5
R1375 VSS.n4916 VSS.n4826 292.5
R1376 VSS.n4929 VSS.n4928 292.5
R1377 VSS.n4932 VSS.n4931 292.5
R1378 VSS.n662 VSS.n661 292.5
R1379 VSS.n659 VSS.n658 292.5
R1380 VSS.n1917 VSS.n1916 292.5
R1381 VSS.n1106 VSS.n147 292.5
R1382 VSS.n1104 VSS.n1103 292.5
R1383 VSS.n1073 VSS.n1072 292.5
R1384 VSS.n1092 VSS.n1091 292.5
R1385 VSS.n1089 VSS.n1088 292.5
R1386 VSS.n1083 VSS.n1082 292.5
R1387 VSS.n1064 VSS.n1058 292.5
R1388 VSS.n4147 VSS.n1057 292.5
R1389 VSS.n4150 VSS.n4149 292.5
R1390 VSS.n4142 VSS.n4141 292.5
R1391 VSS.n4255 VSS.n4254 292.5
R1392 VSS.n4310 VSS.n4309 292.5
R1393 VSS.n4305 VSS.n4304 292.5
R1394 VSS.n4261 VSS.n4260 292.5
R1395 VSS.n4268 VSS.n4262 292.5
R1396 VSS.n4271 VSS.n4264 292.5
R1397 VSS.n4270 VSS.n4263 292.5
R1398 VSS.n4277 VSS.n4265 292.5
R1399 VSS.n4280 VSS.n4279 292.5
R1400 VSS.n4274 VSS.n1040 292.5
R1401 VSS.n4273 VSS.n1039 292.5
R1402 VSS.n4119 VSS.n32 292.5
R1403 VSS.n3055 VSS.n3054 292.5
R1404 VSS.n3054 VSS.n3053 292.5
R1405 VSS.n1459 VSS.n1457 292.5
R1406 VSS.n3052 VSS.n1459 292.5
R1407 VSS.n3050 VSS.n3049 292.5
R1408 VSS.n3051 VSS.n3050 292.5
R1409 VSS.n3021 VSS.n1462 292.5
R1410 VSS.n1462 VSS.n1461 292.5
R1411 VSS.n3004 VSS.n3003 292.5
R1412 VSS.n3003 VSS.n3002 292.5
R1413 VSS.n3000 VSS.n2997 292.5
R1414 VSS.n3001 VSS.n2997 292.5
R1415 VSS.n3032 VSS.n3031 292.5
R1416 VSS.n3033 VSS.n3032 292.5
R1417 VSS.n3008 VSS.n2992 292.5
R1418 VSS.n3034 VSS.n2992 292.5
R1419 VSS.n3037 VSS.n3036 292.5
R1420 VSS.n3036 VSS.n3035 292.5
R1421 VSS.n2991 VSS.n1486 292.5
R1422 VSS.n2996 VSS.n2991 292.5
R1423 VSS.n2994 VSS.n1485 292.5
R1424 VSS.n2993 VSS.n294 292.5
R1425 VSS.n2469 VSS.n2468 292.5
R1426 VSS.n2472 VSS.n2471 292.5
R1427 VSS.n2474 VSS.n1697 292.5
R1428 VSS.n2477 VSS.n2476 292.5
R1429 VSS.n1693 VSS.n1692 292.5
R1430 VSS.n1689 VSS.n1592 292.5
R1431 VSS.n1687 VSS.n1591 292.5
R1432 VSS.n2492 VSS.n2491 292.5
R1433 VSS.n2495 VSS.n2494 292.5
R1434 VSS.n1683 VSS.n1578 292.5
R1435 VSS.n1685 VSS.n1577 292.5
R1436 VSS.n1682 VSS.n1681 292.5
R1437 VSS.n364 VSS.n362 292.5
R1438 VSS.n2360 VSS.n2359 292.5
R1439 VSS.n2355 VSS.n2354 292.5
R1440 VSS.n2106 VSS.n2075 292.5
R1441 VSS.n2100 VSS.n2099 292.5
R1442 VSS.n2091 VSS.n2090 292.5
R1443 VSS.n2088 VSS.n2087 292.5
R1444 VSS.n2072 VSS.n2011 292.5
R1445 VSS.n2070 VSS.n2010 292.5
R1446 VSS.n2460 VSS.n2459 292.5
R1447 VSS.n2463 VSS.n2462 292.5
R1448 VSS.n2466 VSS.n2465 292.5
R1449 VSS.n5366 VSS.n5365 292.5
R1450 VSS.n325 VSS.n324 292.5
R1451 VSS.n5317 VSS.n5316 292.5
R1452 VSS.n2687 VSS.n322 292.5
R1453 VSS.n2693 VSS.n2692 292.5
R1454 VSS.n2683 VSS.n2682 292.5
R1455 VSS.n5322 VSS.n5321 292.5
R1456 VSS.n316 VSS.n312 292.5
R1457 VSS.n319 VSS.n311 292.5
R1458 VSS.n318 VSS.n317 292.5
R1459 VSS.n5360 VSS.n5359 292.5
R1460 VSS.n5363 VSS.n5362 292.5
R1461 VSS.n2726 VSS.n2725 292.5
R1462 VSS.n2721 VSS.n2720 292.5
R1463 VSS.n2669 VSS.n2643 292.5
R1464 VSS.n2664 VSS.n2663 292.5
R1465 VSS.n2655 VSS.n2654 292.5
R1466 VSS.n2653 VSS.n2652 292.5
R1467 VSS.n2640 VSS.n169 292.5
R1468 VSS.n168 VSS.n167 292.5
R1469 VSS.n5423 VSS.n5422 292.5
R1470 VSS.n163 VSS.n159 292.5
R1471 VSS.n5376 VSS.n5375 292.5
R1472 VSS.n5379 VSS.n5378 292.5
R1473 VSS.n5382 VSS.n5381 292.5
R1474 VSS.n5389 VSS.n5388 292.5
R1475 VSS.n5392 VSS.n5391 292.5
R1476 VSS.n229 VSS.n228 292.5
R1477 VSS.n221 VSS.n201 292.5
R1478 VSS.n5403 VSS.n5402 292.5
R1479 VSS.n5406 VSS.n5405 292.5
R1480 VSS.n3343 VSS.n192 292.5
R1481 VSS.n3345 VSS.n191 292.5
R1482 VSS.n3348 VSS.n3347 292.5
R1483 VSS.n3839 VSS.n3838 292.5
R1484 VSS.n3392 VSS.n3391 292.5
R1485 VSS.n3395 VSS.n3394 292.5
R1486 VSS.n3384 VSS.n3383 292.5
R1487 VSS.n3381 VSS.n3380 292.5
R1488 VSS.n3408 VSS.n3407 292.5
R1489 VSS.n3411 VSS.n3410 292.5
R1490 VSS.n3372 VSS.n3371 292.5
R1491 VSS.n3369 VSS.n3368 292.5
R1492 VSS.n3505 VSS.n3504 292.5
R1493 VSS.n1305 VSS.n1304 292.5
R1494 VSS.n3871 VSS.n3870 292.5
R1495 VSS.n1315 VSS.n1310 292.5
R1496 VSS.n3866 VSS.n3865 292.5
R1497 VSS.n3457 VSS.n1313 292.5
R1498 VSS.n3455 VSS.n3454 292.5
R1499 VSS.n3451 VSS.n3450 292.5
R1500 VSS.n3473 VSS.n3472 292.5
R1501 VSS.n3423 VSS.n3422 292.5
R1502 VSS.n3421 VSS.n3420 292.5
R1503 VSS.n1267 VSS.n1266 292.5
R1504 VSS.n1264 VSS.n1263 292.5
R1505 VSS.n1261 VSS.n1260 292.5
R1506 VSS.n1259 VSS.n1258 292.5
R1507 VSS.n1256 VSS.n1255 292.5
R1508 VSS.n1254 VSS.n1253 292.5
R1509 VSS.n1251 VSS.n1250 292.5
R1510 VSS.n1249 VSS.n1248 292.5
R1511 VSS.n1246 VSS.n1245 292.5
R1512 VSS.n996 VSS.n961 292.5
R1513 VSS.n4402 VSS.n4401 292.5
R1514 VSS.n3802 VSS.n1003 292.5
R1515 VSS.n3805 VSS.n3804 292.5
R1516 VSS.n3807 VSS.n3806 292.5
R1517 VSS.n3810 VSS.n3809 292.5
R1518 VSS.n3812 VSS.n3811 292.5
R1519 VSS.n3815 VSS.n3814 292.5
R1520 VSS.n3817 VSS.n3816 292.5
R1521 VSS.n3820 VSS.n3819 292.5
R1522 VSS.n3822 VSS.n3821 292.5
R1523 VSS.n3825 VSS.n3824 292.5
R1524 VSS.n3827 VSS.n3826 292.5
R1525 VSS.n3830 VSS.n3829 292.5
R1526 VSS.n3832 VSS.n3831 292.5
R1527 VSS.n3282 VSS.n3281 292.5
R1528 VSS.n3284 VSS.n3283 292.5
R1529 VSS.n3287 VSS.n3286 292.5
R1530 VSS.n3289 VSS.n3288 292.5
R1531 VSS.n3292 VSS.n3291 292.5
R1532 VSS.n3294 VSS.n3293 292.5
R1533 VSS.n3297 VSS.n3296 292.5
R1534 VSS.n3299 VSS.n3298 292.5
R1535 VSS.n3302 VSS.n3301 292.5
R1536 VSS.n3304 VSS.n3303 292.5
R1537 VSS.n3307 VSS.n3306 292.5
R1538 VSS.n3332 VSS.n3331 292.5
R1539 VSS.n3329 VSS.n3328 292.5
R1540 VSS.n3327 VSS.n3326 292.5
R1541 VSS.n3324 VSS.n3323 292.5
R1542 VSS.n3322 VSS.n3321 292.5
R1543 VSS.n3319 VSS.n3318 292.5
R1544 VSS.n3317 VSS.n3316 292.5
R1545 VSS.n3314 VSS.n3313 292.5
R1546 VSS.n3312 VSS.n3311 292.5
R1547 VSS.n3309 VSS.n3308 292.5
R1548 VSS.n1007 VSS.n151 292.5
R1549 VSS.n4226 VSS.n4225 292.5
R1550 VSS.n4228 VSS.n4227 292.5
R1551 VSS.n4231 VSS.n4230 292.5
R1552 VSS.n4233 VSS.n4232 292.5
R1553 VSS.n4236 VSS.n4235 292.5
R1554 VSS.n4238 VSS.n4237 292.5
R1555 VSS.n4241 VSS.n4240 292.5
R1556 VSS.n4243 VSS.n4242 292.5
R1557 VSS.n4246 VSS.n4245 292.5
R1558 VSS.n4248 VSS.n4247 292.5
R1559 VSS.n4251 VSS.n4250 292.5
R1560 VSS.n4224 VSS.n4223 292.5
R1561 VSS.n4221 VSS.n4220 292.5
R1562 VSS.n4219 VSS.n4218 292.5
R1563 VSS.n4216 VSS.n4215 292.5
R1564 VSS.n4214 VSS.n4213 292.5
R1565 VSS.n4211 VSS.n4210 292.5
R1566 VSS.n4209 VSS.n4208 292.5
R1567 VSS.n4206 VSS.n4205 292.5
R1568 VSS.n1012 VSS.n1011 292.5
R1569 VSS.n20 VSS.t64 284.349
R1570 VSS.n1 VSS.t61 284.334
R1571 VSS.t36 VSS.n339 284.014
R1572 VSS.n4143 VSS.n1063 272.089
R1573 VSS.n717 VSS.n674 272.089
R1574 VSS.n4665 VSS.n674 272.089
R1575 VSS.n714 VSS.n674 272.089
R1576 VSS.n4674 VSS.n674 272.089
R1577 VSS.n711 VSS.n674 272.089
R1578 VSS.n1896 VSS.n674 272.089
R1579 VSS.n1886 VSS.n674 272.089
R1580 VSS.n1905 VSS.n674 272.089
R1581 VSS.n1883 VSS.n674 272.089
R1582 VSS.n1914 VSS.n674 272.089
R1583 VSS.n1948 VSS.n674 272.089
R1584 VSS.n1943 VSS.n674 272.089
R1585 VSS.n1922 VSS.n674 272.089
R1586 VSS.n1934 VSS.n674 272.089
R1587 VSS.n1929 VSS.n674 272.089
R1588 VSS.n2172 VSS.n674 272.089
R1589 VSS.n2185 VSS.n674 272.089
R1590 VSS.n2169 VSS.n674 272.089
R1591 VSS.n2194 VSS.n674 272.089
R1592 VSS.n2167 VSS.n674 272.089
R1593 VSS.n2202 VSS.n674 272.089
R1594 VSS.n2159 VSS.n674 272.089
R1595 VSS.n2211 VSS.n674 272.089
R1596 VSS.n2156 VSS.n674 272.089
R1597 VSS.n2220 VSS.n674 272.089
R1598 VSS.n2292 VSS.n2291 272.089
R1599 VSS.n4658 VSS.n710 272.089
R1600 VSS.n4663 VSS.n710 272.089
R1601 VSS.n4667 VSS.n710 272.089
R1602 VSS.n4672 VSS.n710 272.089
R1603 VSS.n4676 VSS.n710 272.089
R1604 VSS.n1894 VSS.n710 272.089
R1605 VSS.n1898 VSS.n710 272.089
R1606 VSS.n1903 VSS.n710 272.089
R1607 VSS.n1907 VSS.n710 272.089
R1608 VSS.n1912 VSS.n710 272.089
R1609 VSS.n1950 VSS.n710 272.089
R1610 VSS.n1920 VSS.n710 272.089
R1611 VSS.n1941 VSS.n710 272.089
R1612 VSS.n1936 VSS.n710 272.089
R1613 VSS.n1924 VSS.n710 272.089
R1614 VSS.n2178 VSS.n710 272.089
R1615 VSS.n2183 VSS.n710 272.089
R1616 VSS.n2187 VSS.n710 272.089
R1617 VSS.n2192 VSS.n710 272.089
R1618 VSS.n2196 VSS.n710 272.089
R1619 VSS.n2163 VSS.n710 272.089
R1620 VSS.n2204 VSS.n710 272.089
R1621 VSS.n2209 VSS.n710 272.089
R1622 VSS.n2213 VSS.n710 272.089
R1623 VSS.n2218 VSS.n710 272.089
R1624 VSS.n382 VSS.n374 272.089
R1625 VSS.n5229 VSS.n384 272.089
R1626 VSS.n2402 VSS.n374 272.089
R1627 VSS.n5229 VSS.n385 272.089
R1628 VSS.n2053 VSS.n374 272.089
R1629 VSS.n5229 VSS.n386 272.089
R1630 VSS.n2417 VSS.n374 272.089
R1631 VSS.n5229 VSS.n387 272.089
R1632 VSS.n2040 VSS.n374 272.089
R1633 VSS.n5229 VSS.n388 272.089
R1634 VSS.n390 VSS.n374 272.089
R1635 VSS.n2176 VSS.n674 272.089
R1636 VSS.n1927 VSS.n710 272.089
R1637 VSS.n1795 VSS.n394 272.089
R1638 VSS.n5225 VSS.n395 272.089
R1639 VSS.n1797 VSS.n1795 272.089
R1640 VSS.n5225 VSS.n396 272.089
R1641 VSS.n1795 VSS.n1794 272.089
R1642 VSS.n5225 VSS.n397 272.089
R1643 VSS.n1795 VSS.n1713 272.089
R1644 VSS.n5225 VSS.n398 272.089
R1645 VSS.n1795 VSS.n1712 272.089
R1646 VSS.n5225 VSS.n399 272.089
R1647 VSS.n1795 VSS.n401 272.089
R1648 VSS.n3223 VSS.n1353 272.089
R1649 VSS.n3150 VSS.n3149 272.089
R1650 VSS.n3223 VSS.n1352 272.089
R1651 VSS.n3149 VSS.n3148 272.089
R1652 VSS.n3223 VSS.n1351 272.089
R1653 VSS.n3149 VSS.n1409 272.089
R1654 VSS.n3223 VSS.n1350 272.089
R1655 VSS.n3149 VSS.n1408 272.089
R1656 VSS.n3223 VSS.n1349 272.089
R1657 VSS.n3149 VSS.n1348 272.089
R1658 VSS.n4556 VSS.n4555 272.089
R1659 VSS.n4557 VSS.n792 272.089
R1660 VSS.n835 VSS.n792 272.089
R1661 VSS.n4555 VSS.n805 272.089
R1662 VSS.n4570 VSS.n792 272.089
R1663 VSS.n4555 VSS.n804 272.089
R1664 VSS.n802 VSS.n792 272.089
R1665 VSS.n4555 VSS.n793 272.089
R1666 VSS.n4583 VSS.n792 272.089
R1667 VSS.n4555 VSS.n791 272.089
R1668 VSS.n4553 VSS.n792 272.089
R1669 VSS.n3919 VSS.n244 272.089
R1670 VSS.n3914 VSS.n244 272.089
R1671 VSS.n3909 VSS.n244 272.089
R1672 VSS.n3904 VSS.n244 272.089
R1673 VSS.n3899 VSS.n244 272.089
R1674 VSS.n3226 VSS.n244 272.089
R1675 VSS.n3231 VSS.n244 272.089
R1676 VSS.n3236 VSS.n244 272.089
R1677 VSS.n3241 VSS.n244 272.089
R1678 VSS.n3246 VSS.n244 272.089
R1679 VSS.n3251 VSS.n244 272.089
R1680 VSS.n2871 VSS.n244 272.089
R1681 VSS.n2876 VSS.n244 272.089
R1682 VSS.n2881 VSS.n244 272.089
R1683 VSS.n2886 VSS.n244 272.089
R1684 VSS.n2891 VSS.n244 272.089
R1685 VSS.n2894 VSS.n244 272.089
R1686 VSS.n2900 VSS.n244 272.089
R1687 VSS.n2905 VSS.n244 272.089
R1688 VSS.n2910 VSS.n244 272.089
R1689 VSS.n2915 VSS.n244 272.089
R1690 VSS.n2920 VSS.n244 272.089
R1691 VSS.n2617 VSS.n244 272.089
R1692 VSS.n2614 VSS.n244 272.089
R1693 VSS.n2609 VSS.n244 272.089
R1694 VSS.n2604 VSS.n244 272.089
R1695 VSS.n2599 VSS.n244 272.089
R1696 VSS.n2594 VSS.n244 272.089
R1697 VSS.n1496 VSS.n244 272.089
R1698 VSS.n1501 VSS.n244 272.089
R1699 VSS.n1506 VSS.n244 272.089
R1700 VSS.n1511 VSS.n244 272.089
R1701 VSS.n1514 VSS.n244 272.089
R1702 VSS.n1519 VSS.n1518 272.089
R1703 VSS.n5372 VSS.n272 272.089
R1704 VSS.n5372 VSS.n271 272.089
R1705 VSS.n5372 VSS.n270 272.089
R1706 VSS.n5372 VSS.n269 272.089
R1707 VSS.n5372 VSS.n268 272.089
R1708 VSS.n5372 VSS.n267 272.089
R1709 VSS.n5372 VSS.n273 272.089
R1710 VSS.n5372 VSS.n274 272.089
R1711 VSS.n5372 VSS.n275 272.089
R1712 VSS.n5372 VSS.n276 272.089
R1713 VSS.n5372 VSS.n277 272.089
R1714 VSS.n5372 VSS.n278 272.089
R1715 VSS.n5372 VSS.n265 272.089
R1716 VSS.n5372 VSS.n264 272.089
R1717 VSS.n5372 VSS.n263 272.089
R1718 VSS.n5372 VSS.n262 272.089
R1719 VSS.n5372 VSS.n261 272.089
R1720 VSS.n5372 VSS.n260 272.089
R1721 VSS.n5372 VSS.n280 272.089
R1722 VSS.n5372 VSS.n281 272.089
R1723 VSS.n5372 VSS.n282 272.089
R1724 VSS.n5372 VSS.n283 272.089
R1725 VSS.n5372 VSS.n284 272.089
R1726 VSS.n5372 VSS.n257 272.089
R1727 VSS.n5372 VSS.n256 272.089
R1728 VSS.n5372 VSS.n255 272.089
R1729 VSS.n5372 VSS.n254 272.089
R1730 VSS.n5372 VSS.n253 272.089
R1731 VSS.n5372 VSS.n252 272.089
R1732 VSS.n5372 VSS.n286 272.089
R1733 VSS.n5372 VSS.n287 272.089
R1734 VSS.n5372 VSS.n288 272.089
R1735 VSS.n5372 VSS.n289 272.089
R1736 VSS.n4464 VSS.n406 272.089
R1737 VSS.n4488 VSS.n406 272.089
R1738 VSS.n4483 VSS.n406 272.089
R1739 VSS.n4468 VSS.n406 272.089
R1740 VSS.n4474 VSS.n406 272.089
R1741 VSS.n3187 VSS.n406 272.089
R1742 VSS.n3194 VSS.n406 272.089
R1743 VSS.n3184 VSS.n406 272.089
R1744 VSS.n3203 VSS.n406 272.089
R1745 VSS.n3181 VSS.n406 272.089
R1746 VSS.n3212 VSS.n406 272.089
R1747 VSS.n5200 VSS.n406 272.089
R1748 VSS.n412 VSS.n406 272.089
R1749 VSS.n5209 VSS.n406 272.089
R1750 VSS.n409 VSS.n406 272.089
R1751 VSS.n5218 VSS.n406 272.089
R1752 VSS.n1622 VSS.n406 272.089
R1753 VSS.n1629 VSS.n406 272.089
R1754 VSS.n1619 VSS.n406 272.089
R1755 VSS.n1638 VSS.n406 272.089
R1756 VSS.n1616 VSS.n406 272.089
R1757 VSS.n1647 VSS.n406 272.089
R1758 VSS.n1652 VSS.n406 272.089
R1759 VSS.n1671 VSS.n406 272.089
R1760 VSS.n1666 VSS.n406 272.089
R1761 VSS.n1656 VSS.n406 272.089
R1762 VSS.n1657 VSS.n406 272.089
R1763 VSS.n2533 VSS.n1559 272.089
R1764 VSS.n4496 VSS.n407 272.089
R1765 VSS.n4490 VSS.n407 272.089
R1766 VSS.n4466 VSS.n407 272.089
R1767 VSS.n4481 VSS.n407 272.089
R1768 VSS.n4476 VSS.n407 272.089
R1769 VSS.n4471 VSS.n407 272.089
R1770 VSS.n3192 VSS.n407 272.089
R1771 VSS.n3196 VSS.n407 272.089
R1772 VSS.n3201 VSS.n407 272.089
R1773 VSS.n3205 VSS.n407 272.089
R1774 VSS.n3210 VSS.n407 272.089
R1775 VSS.n3214 VSS.n407 272.089
R1776 VSS.n414 VSS.n407 272.089
R1777 VSS.n5202 VSS.n407 272.089
R1778 VSS.n5207 VSS.n407 272.089
R1779 VSS.n5211 VSS.n407 272.089
R1780 VSS.n5216 VSS.n407 272.089
R1781 VSS.n5220 VSS.n407 272.089
R1782 VSS.n1627 VSS.n407 272.089
R1783 VSS.n1631 VSS.n407 272.089
R1784 VSS.n1636 VSS.n407 272.089
R1785 VSS.n1640 VSS.n407 272.089
R1786 VSS.n1645 VSS.n407 272.089
R1787 VSS.n1678 VSS.n407 272.089
R1788 VSS.n1673 VSS.n407 272.089
R1789 VSS.n1654 VSS.n407 272.089
R1790 VSS.n1664 VSS.n407 272.089
R1791 VSS.n1659 VSS.n407 272.089
R1792 VSS.n1383 VSS.n406 272.089
R1793 VSS.n1358 VSS.n406 272.089
R1794 VSS.n1374 VSS.n406 272.089
R1795 VSS.n1369 VSS.n406 272.089
R1796 VSS.n1364 VSS.n406 272.089
R1797 VSS.n1381 VSS.n407 272.089
R1798 VSS.n1376 VSS.n407 272.089
R1799 VSS.n1360 VSS.n407 272.089
R1800 VSS.n1367 VSS.n407 272.089
R1801 VSS.n1362 VSS.n407 272.089
R1802 VSS.n3149 VSS.n1354 272.089
R1803 VSS.n1356 VSS.n407 272.089
R1804 VSS.n497 VSS.n454 272.089
R1805 VSS.n5124 VSS.n456 272.089
R1806 VSS.n492 VSS.n456 272.089
R1807 VSS.n490 VSS.n454 272.089
R1808 VSS.n488 VSS.n456 272.089
R1809 VSS.n457 VSS.n454 272.089
R1810 VSS.n5148 VSS.n456 272.089
R1811 VSS.n5150 VSS.n454 272.089
R1812 VSS.n456 VSS.n453 272.089
R1813 VSS.n3219 VSS.n454 272.089
R1814 VSS.n4878 VSS.n621 272.089
R1815 VSS.n5120 VSS.n504 272.089
R1816 VSS.n4870 VSS.n621 272.089
R1817 VSS.n5120 VSS.n505 272.089
R1818 VSS.n4861 VSS.n621 272.089
R1819 VSS.n5120 VSS.n506 272.089
R1820 VSS.n4848 VSS.n621 272.089
R1821 VSS.n5120 VSS.n507 272.089
R1822 VSS.n621 VSS.n509 272.089
R1823 VSS.n5120 VSS.n5119 272.089
R1824 VSS.n621 VSS.n502 272.089
R1825 VSS.n1889 VSS.n674 272.089
R1826 VSS.n684 VSS.n674 272.089
R1827 VSS.n700 VSS.n674 272.089
R1828 VSS.n695 VSS.n674 272.089
R1829 VSS.n690 VSS.n674 272.089
R1830 VSS.n680 VSS.n674 272.089
R1831 VSS.n710 VSS.n709 272.089
R1832 VSS.n710 VSS.n679 272.089
R1833 VSS.n710 VSS.n678 272.089
R1834 VSS.n710 VSS.n677 272.089
R1835 VSS.n710 VSS.n676 272.089
R1836 VSS.n682 VSS.n674 272.089
R1837 VSS.n4681 VSS.n710 272.089
R1838 VSS.n4740 VSS.n4691 272.089
R1839 VSS.n4779 VSS.n4778 272.089
R1840 VSS.n4740 VSS.n4733 272.089
R1841 VSS.n4779 VSS.n4689 272.089
R1842 VSS.n4740 VSS.n4736 272.089
R1843 VSS.n4779 VSS.n4688 272.089
R1844 VSS.n4740 VSS.n4739 272.089
R1845 VSS.n4779 VSS.n4687 272.089
R1846 VSS.n4741 VSS.n4740 272.089
R1847 VSS.n4779 VSS.n4686 272.089
R1848 VSS.n4740 VSS.n4684 272.089
R1849 VSS.n3923 VSS.n3896 272.089
R1850 VSS.n4498 VSS.n4463 272.089
R1851 VSS.n736 VSS.n719 272.089
R1852 VSS.n1269 VSS.n1243 272.089
R1853 VSS.n3758 VSS.n3582 272.089
R1854 VSS.n3708 VSS.n3582 272.089
R1855 VSS.n3710 VSS.n3587 272.089
R1856 VSS.n3673 VSS.n3582 272.089
R1857 VSS.n3710 VSS.n3586 272.089
R1858 VSS.n3664 VSS.n3582 272.089
R1859 VSS.n3710 VSS.n3585 272.089
R1860 VSS.n3655 VSS.n3582 272.089
R1861 VSS.n3710 VSS.n3581 272.089
R1862 VSS.n3710 VSS.n3584 272.089
R1863 VSS.n3797 VSS.n3796 272.089
R1864 VSS.n4020 VSS.n1122 272.089
R1865 VSS.n3796 VSS.n3524 272.089
R1866 VSS.n4020 VSS.n1121 272.089
R1867 VSS.n3796 VSS.n3525 272.089
R1868 VSS.n4020 VSS.n1120 272.089
R1869 VSS.n3796 VSS.n3526 272.089
R1870 VSS.n4020 VSS.n1119 272.089
R1871 VSS.n3796 VSS.n3795 272.089
R1872 VSS.n4021 VSS.n4020 272.089
R1873 VSS.n3796 VSS.n1117 272.089
R1874 VSS.n5456 VSS.n5455 272.089
R1875 VSS.n5473 VSS.n78 272.089
R1876 VSS.n5455 VSS.n5454 272.089
R1877 VSS.n5473 VSS.n79 272.089
R1878 VSS.n5455 VSS.n116 272.089
R1879 VSS.n5473 VSS.n80 272.089
R1880 VSS.n5455 VSS.n115 272.089
R1881 VSS.n5473 VSS.n81 272.089
R1882 VSS.n5455 VSS.n83 272.089
R1883 VSS.n5473 VSS.n5472 272.089
R1884 VSS.n5455 VSS.n75 272.089
R1885 VSS.n245 VSS.n241 272.089
R1886 VSS.n258 VSS.n241 272.089
R1887 VSS.n5192 VSS.n416 272.089
R1888 VSS.n5194 VSS.n416 272.089
R1889 VSS.n1875 VSS.n1874 272.089
R1890 VSS.n5189 VSS.n423 272.089
R1891 VSS.n1874 VSS.n1873 272.089
R1892 VSS.n5189 VSS.n424 272.089
R1893 VSS.n1874 VSS.n1813 272.089
R1894 VSS.n5189 VSS.n425 272.089
R1895 VSS.n1874 VSS.n1812 272.089
R1896 VSS.n5189 VSS.n426 272.089
R1897 VSS.n1874 VSS.n428 272.089
R1898 VSS.n5189 VSS.n5188 272.089
R1899 VSS.n1874 VSS.n421 272.089
R1900 VSS.n1954 VSS.n1879 272.089
R1901 VSS.n1954 VSS.n1878 272.089
R1902 VSS.n4949 VSS.n4948 272.089
R1903 VSS.n4945 VSS.n620 272.089
R1904 VSS.n4948 VSS.n4947 272.089
R1905 VSS.n4909 VSS.n620 272.089
R1906 VSS.n4948 VSS.n633 272.089
R1907 VSS.n4917 VSS.n620 272.089
R1908 VSS.n4948 VSS.n632 272.089
R1909 VSS.n4930 VSS.n620 272.089
R1910 VSS.n4948 VSS.n631 272.089
R1911 VSS.n660 VSS.n620 272.089
R1912 VSS.n4948 VSS.n630 272.089
R1913 VSS.n1105 VSS.n1063 272.089
R1914 VSS.n4145 VSS.n1107 272.089
R1915 VSS.n1067 VSS.n1063 272.089
R1916 VSS.n4145 VSS.n1066 272.089
R1917 VSS.n1090 VSS.n1063 272.089
R1918 VSS.n4145 VSS.n1065 272.089
R1919 VSS.n1081 VSS.n1063 272.089
R1920 VSS.n4146 VSS.n4145 272.089
R1921 VSS.n4148 VSS.n1063 272.089
R1922 VSS.n4145 VSS.n1062 272.089
R1923 VSS.n4308 VSS.n4307 272.089
R1924 VSS.n4276 VSS.n4200 272.089
R1925 VSS.n4307 VSS.n4306 272.089
R1926 VSS.n4276 VSS.n4269 272.089
R1927 VSS.n4307 VSS.n4259 272.089
R1928 VSS.n4276 VSS.n4272 272.089
R1929 VSS.n4307 VSS.n4258 272.089
R1930 VSS.n4278 VSS.n4276 272.089
R1931 VSS.n4307 VSS.n4257 272.089
R1932 VSS.n4276 VSS.n4275 272.089
R1933 VSS.n4307 VSS.n4256 272.089
R1934 VSS.n5367 VSS.n292 272.089
R1935 VSS.n5368 VSS.n5367 272.089
R1936 VSS.n1649 VSS.n1458 272.089
R1937 VSS.n1651 VSS.n1458 272.089
R1938 VSS.n1698 VSS.n1695 272.089
R1939 VSS.n2473 VSS.n1584 272.089
R1940 VSS.n2475 VSS.n1695 272.089
R1941 VSS.n1612 VSS.n1584 272.089
R1942 VSS.n1695 VSS.n1694 272.089
R1943 VSS.n1688 VSS.n1584 272.089
R1944 VSS.n1695 VSS.n1585 272.089
R1945 VSS.n2493 VSS.n1584 272.089
R1946 VSS.n1695 VSS.n1583 272.089
R1947 VSS.n1684 VSS.n1584 272.089
R1948 VSS.n1695 VSS.n1686 272.089
R1949 VSS.n2165 VSS.n1997 272.089
R1950 VSS.n2161 VSS.n1997 272.089
R1951 VSS.n2358 VSS.n2357 272.089
R1952 VSS.n2069 VSS.n373 272.089
R1953 VSS.n2357 VSS.n2356 272.089
R1954 VSS.n2098 VSS.n373 272.089
R1955 VSS.n2357 VSS.n2074 272.089
R1956 VSS.n2089 VSS.n373 272.089
R1957 VSS.n2357 VSS.n2073 272.089
R1958 VSS.n2071 VSS.n373 272.089
R1959 VSS.n2357 VSS.n2005 272.089
R1960 VSS.n2461 VSS.n373 272.089
R1961 VSS.n2357 VSS.n2000 272.089
R1962 VSS.n5319 VSS.n296 272.089
R1963 VSS.n5364 VSS.n297 272.089
R1964 VSS.n5319 VSS.n5318 272.089
R1965 VSS.n5364 VSS.n298 272.089
R1966 VSS.n5319 VSS.n321 272.089
R1967 VSS.n5364 VSS.n299 272.089
R1968 VSS.n5320 VSS.n5319 272.089
R1969 VSS.n5364 VSS.n300 272.089
R1970 VSS.n5319 VSS.n320 272.089
R1971 VSS.n5364 VSS.n301 272.089
R1972 VSS.n5319 VSS.n303 272.089
R1973 VSS.n2724 VSS.n2723 272.089
R1974 VSS.n5425 VSS.n155 272.089
R1975 VSS.n2723 VSS.n2722 272.089
R1976 VSS.n5425 VSS.n156 272.089
R1977 VSS.n2723 VSS.n2642 272.089
R1978 VSS.n5425 VSS.n157 272.089
R1979 VSS.n2723 VSS.n2641 272.089
R1980 VSS.n5425 VSS.n158 272.089
R1981 VSS.n2723 VSS.n160 272.089
R1982 VSS.n5425 VSS.n5424 272.089
R1983 VSS.n2723 VSS.n153 272.089
R1984 VSS.n3342 VSS.n234 272.089
R1985 VSS.n5380 VSS.n198 272.089
R1986 VSS.n3342 VSS.n231 272.089
R1987 VSS.n5390 VSS.n198 272.089
R1988 VSS.n3342 VSS.n230 272.089
R1989 VSS.n222 VSS.n198 272.089
R1990 VSS.n3342 VSS.n199 272.089
R1991 VSS.n5404 VSS.n198 272.089
R1992 VSS.n3342 VSS.n197 272.089
R1993 VSS.n3344 VSS.n198 272.089
R1994 VSS.n3346 VSS.n3342 272.089
R1995 VSS.n3837 VSS.n1344 272.089
R1996 VSS.n3835 VSS.n1343 272.089
R1997 VSS.n3393 VSS.n1344 272.089
R1998 VSS.n3835 VSS.n3257 272.089
R1999 VSS.n3382 VSS.n1344 272.089
R2000 VSS.n3835 VSS.n3258 272.089
R2001 VSS.n3409 VSS.n1344 272.089
R2002 VSS.n3835 VSS.n3259 272.089
R2003 VSS.n3370 VSS.n1344 272.089
R2004 VSS.n3835 VSS.n3260 272.089
R2005 VSS.n3262 VSS.n1344 272.089
R2006 VSS.n3868 VSS.n948 272.089
R2007 VSS.n4405 VSS.n951 272.089
R2008 VSS.n3869 VSS.n3868 272.089
R2009 VSS.n4405 VSS.n952 272.089
R2010 VSS.n3868 VSS.n3867 272.089
R2011 VSS.n4405 VSS.n953 272.089
R2012 VSS.n3868 VSS.n1312 272.089
R2013 VSS.n4405 VSS.n954 272.089
R2014 VSS.n3868 VSS.n1311 272.089
R2015 VSS.n4405 VSS.n955 272.089
R2016 VSS.n3868 VSS.n957 272.089
R2017 VSS.n1265 VSS.n1008 272.089
R2018 VSS.n1262 VSS.n1008 272.089
R2019 VSS.n1257 VSS.n1008 272.089
R2020 VSS.n1252 VSS.n1008 272.089
R2021 VSS.n1247 VSS.n1008 272.089
R2022 VSS.n1008 VSS.n962 272.089
R2023 VSS.n3803 VSS.n1008 272.089
R2024 VSS.n3808 VSS.n1008 272.089
R2025 VSS.n3813 VSS.n1008 272.089
R2026 VSS.n3818 VSS.n1008 272.089
R2027 VSS.n3823 VSS.n1008 272.089
R2028 VSS.n3828 VSS.n1008 272.089
R2029 VSS.n3285 VSS.n1008 272.089
R2030 VSS.n3290 VSS.n1008 272.089
R2031 VSS.n3295 VSS.n1008 272.089
R2032 VSS.n3300 VSS.n1008 272.089
R2033 VSS.n3305 VSS.n1008 272.089
R2034 VSS.n3337 VSS.n3336 272.089
R2035 VSS.n3338 VSS.n3337 272.089
R2036 VSS.n3330 VSS.n1008 272.089
R2037 VSS.n3325 VSS.n1008 272.089
R2038 VSS.n3320 VSS.n1008 272.089
R2039 VSS.n3315 VSS.n1008 272.089
R2040 VSS.n3310 VSS.n1008 272.089
R2041 VSS.n4229 VSS.n1008 272.089
R2042 VSS.n4234 VSS.n1008 272.089
R2043 VSS.n4239 VSS.n1008 272.089
R2044 VSS.n4244 VSS.n1008 272.089
R2045 VSS.n4249 VSS.n1008 272.089
R2046 VSS.n4253 VSS.n4204 272.089
R2047 VSS.n4253 VSS.n4202 272.089
R2048 VSS.n4222 VSS.n1008 272.089
R2049 VSS.n4217 VSS.n1008 272.089
R2050 VSS.n4212 VSS.n1008 272.089
R2051 VSS.n4207 VSS.n1008 272.089
R2052 VSS.n4330 VSS.n1009 272.089
R2053 VSS.n1010 VSS.n1008 272.089
R2054 VSS.n4400 VSS.n1001 272.089
R2055 VSS.n4400 VSS.n1000 272.089
R2056 VSS.n4400 VSS.n999 272.089
R2057 VSS.n4400 VSS.n998 272.089
R2058 VSS.n4400 VSS.n997 272.089
R2059 VSS.n4400 VSS.n995 272.089
R2060 VSS.n4400 VSS.n994 272.089
R2061 VSS.n4400 VSS.n993 272.089
R2062 VSS.n4400 VSS.n992 272.089
R2063 VSS.n4400 VSS.n991 272.089
R2064 VSS.n4400 VSS.n990 272.089
R2065 VSS.n4400 VSS.n989 272.089
R2066 VSS.n4400 VSS.n988 272.089
R2067 VSS.n4400 VSS.n987 272.089
R2068 VSS.n4400 VSS.n986 272.089
R2069 VSS.n4400 VSS.n985 272.089
R2070 VSS.n4400 VSS.n984 272.089
R2071 VSS.n4400 VSS.n982 272.089
R2072 VSS.n4400 VSS.n981 272.089
R2073 VSS.n4400 VSS.n980 272.089
R2074 VSS.n4400 VSS.n979 272.089
R2075 VSS.n4400 VSS.n978 272.089
R2076 VSS.n4400 VSS.n977 272.089
R2077 VSS.n4400 VSS.n976 272.089
R2078 VSS.n4400 VSS.n975 272.089
R2079 VSS.n4400 VSS.n974 272.089
R2080 VSS.n4400 VSS.n973 272.089
R2081 VSS.n4400 VSS.n972 272.089
R2082 VSS.n4400 VSS.n971 272.089
R2083 VSS.n4400 VSS.n969 272.089
R2084 VSS.n4400 VSS.n968 272.089
R2085 VSS.n4400 VSS.n967 272.089
R2086 VSS.n4400 VSS.n966 272.089
R2087 VSS.n4400 VSS.n965 272.089
R2088 VSS.n1099 VSS.n145 258.334
R2089 VSS.n3549 VSS.n3548 258.334
R2090 VSS.n3703 VSS.n3684 258.334
R2091 VSS.n3876 VSS.n3875 258.334
R2092 VSS.n4898 VSS.n4897 258.334
R2093 VSS.n1866 VSS.n1865 258.334
R2094 VSS.n5128 VSS.n483 258.334
R2095 VSS.n2079 VSS.n2066 258.334
R2096 VSS.n1699 VSS.n1607 258.334
R2097 VSS.n3014 VSS.n1455 258.334
R2098 VSS.n2701 VSS.n2700 258.334
R2099 VSS.n3124 VSS.n3123 258.334
R2100 VSS.n235 VSS.n217 258.334
R2101 VSS.n1183 VSS.t7 257.493
R2102 VSS.n5562 VSS.n6 257.466
R2103 VSS.n5279 VSS.n350 254.34
R2104 VSS.n5014 VSS.n611 254.34
R2105 VSS.n5066 VSS.n583 254.34
R2106 VSS.n3994 VSS.n3993 254.34
R2107 VSS.n1211 VSS.n1202 254.34
R2108 VSS.n1212 VSS.n1211 254.34
R2109 VSS.n1211 VSS.n1210 254.34
R2110 VSS.n4991 VSS.n4990 254.34
R2111 VSS.n5256 VSS.n5255 254.34
R2112 VSS.n1135 VSS.n71 254.34
R2113 VSS.n33 VSS.n28 254.34
R2114 VSS.n5561 VSS.n7 254.34
R2115 VSS.n4315 VSS.n1041 250
R2116 VSS.n4042 VSS.n4041 250
R2117 VSS.n5104 VSS.n540 250
R2118 VSS.n4798 VSS.n4797 250
R2119 VSS.n4588 VSS.n4587 250
R2120 VSS.n4535 VSS.n869 250
R2121 VSS.n2033 VSS.n2032 250
R2122 VSS.n2302 VSS.n2131 250
R2123 VSS.n2519 VSS.n2518 250
R2124 VSS.n2563 VSS.n2562 250
R2125 VSS.n4387 VSS.n4386 250
R2126 VSS.n4104 VSS.n4103 250
R2127 VSS.n1765 VSS.n1763 250
R2128 VSS.n2967 VSS.n2587 250
R2129 VSS.n3266 VSS.n3265 250
R2130 VSS.n2789 VSS.n2788 250
R2131 VSS.n3496 VSS.n3495 250
R2132 VSS.n5280 VSS.n349 249.663
R2133 VSS.n52 VSS.n51 240.334
R2134 VSS.n1177 VSS.t52 228.215
R2135 VSS.n1176 VSS.t51 228.215
R2136 VSS.n1175 VSS.t50 228.215
R2137 VSS.n1174 VSS.t49 228.215
R2138 VSS.t7 VSS.n341 226.368
R2139 VSS.n1101 VSS.n1051 221.667
R2140 VSS.n5447 VSS.n5446 221.667
R2141 VSS.n3562 VSS.n101 221.667
R2142 VSS.n3607 VSS.n3606 221.667
R2143 VSS.n3967 VSS.n1240 221.667
R2144 VSS.n3891 VSS.n1299 221.667
R2145 VSS.n5076 VSS.n5075 221.667
R2146 VSS.n4772 VSS.n4771 221.667
R2147 VSS.n4883 VSS.n4838 221.667
R2148 VSS.n1851 VSS.n1850 221.667
R2149 VSS.n832 VSS.n831 221.667
R2150 VSS.n4642 VSS.n4641 221.667
R2151 VSS.n4507 VSS.n4506 221.667
R2152 VSS.n2398 VSS.n2397 221.667
R2153 VSS.n4942 VSS.n4941 221.667
R2154 VSS.n2352 VSS.n2351 221.667
R2155 VSS.n2264 VSS.n2263 221.667
R2156 VSS.n3047 VSS.n3046 221.667
R2157 VSS.n5314 VSS.n5313 221.667
R2158 VSS.n4197 VSS.n4196 221.667
R2159 VSS.n1980 VSS.n1979 221.667
R2160 VSS.n1958 VSS.n1808 221.667
R2161 VSS.n3074 VSS.n3073 221.667
R2162 VSS.n3106 VSS.n3105 221.667
R2163 VSS.n2718 VSS.n2717 221.667
R2164 VSS.n238 VSS.n237 221.667
R2165 VSS.n3141 VSS.n3140 221.667
R2166 VSS.n4542 VSS.n4541 221.667
R2167 VSS.n1340 VSS.n1339 221.667
R2168 VSS.n3860 VSS.n3859 221.667
R2169 VSS.n4307 VSS.n31 221.278
R2170 VSS.n5455 VSS.n73 221.278
R2171 VSS.n3752 VSS.n3710 221.278
R2172 VSS.n4020 VSS.n1124 221.278
R2173 VSS.n4145 VSS.n59 221.278
R2174 VSS.n4877 VSS.n607 213.333
R2175 VSS.n22 VSS.t94 213.059
R2176 VSS.n4008 VSS.t91 213.042
R2177 VSS.n5288 VSS.n338 210.599
R2178 VSS.n4276 VSS.n31 208.512
R2179 VSS.n5473 VSS.n73 208.512
R2180 VSS.n3752 VSS.n3582 208.512
R2181 VSS.n3796 VSS.n1124 208.512
R2182 VSS.n1063 VSS.n59 208.512
R2183 VSS.n5281 VSS.n348 204.757
R2184 VSS.n5276 VSS.n348 204.757
R2185 VSS.n5276 VSS.n5275 204.757
R2186 VSS.n5275 VSS.n5274 204.757
R2187 VSS.n5274 VSS.n353 204.757
R2188 VSS.n5268 VSS.n5267 204.757
R2189 VSS.n5267 VSS.n5266 204.757
R2190 VSS.n5266 VSS.n358 204.757
R2191 VSS.n5260 VSS.n358 204.757
R2192 VSS.n5260 VSS.n5259 204.757
R2193 VSS.n5259 VSS.n5258 204.757
R2194 VSS.n5253 VSS.n367 204.757
R2195 VSS.n5253 VSS.n5252 204.757
R2196 VSS.n5252 VSS.n5251 204.757
R2197 VSS.n5251 VSS.n368 204.757
R2198 VSS.n5245 VSS.n368 204.757
R2199 VSS.n5244 VSS.n5243 204.757
R2200 VSS.n5243 VSS.n375 204.757
R2201 VSS.n5237 VSS.n375 204.757
R2202 VSS.n5237 VSS.n5236 204.757
R2203 VSS.n5236 VSS.n5235 204.757
R2204 VSS.n5235 VSS.n379 204.757
R2205 VSS.n4965 VSS.n4964 204.757
R2206 VSS.n4965 VSS.n4960 204.757
R2207 VSS.n4972 VSS.n4960 204.757
R2208 VSS.n4973 VSS.n4972 204.757
R2209 VSS.n4974 VSS.n4973 204.757
R2210 VSS.n4978 VSS.n4977 204.757
R2211 VSS.n4978 VSS.n4955 204.757
R2212 VSS.n4985 VSS.n4955 204.757
R2213 VSS.n4986 VSS.n4985 204.757
R2214 VSS.n4988 VSS.n4986 204.757
R2215 VSS.n4988 VSS.n4987 204.757
R2216 VSS.n4993 VSS.n626 204.757
R2217 VSS.n4994 VSS.n4993 204.757
R2218 VSS.n4995 VSS.n4994 204.757
R2219 VSS.n4995 VSS.n622 204.757
R2220 VSS.n5001 VSS.n622 204.757
R2221 VSS.n5003 VSS.n5002 204.757
R2222 VSS.n5003 VSS.n616 204.757
R2223 VSS.n5009 VSS.n616 204.757
R2224 VSS.n5010 VSS.n5009 204.757
R2225 VSS.n5012 VSS.n5010 204.757
R2226 VSS.n5012 VSS.n5011 204.757
R2227 VSS.n613 VSS.n605 204.757
R2228 VSS.n5019 VSS.n605 204.757
R2229 VSS.n5020 VSS.n5019 204.757
R2230 VSS.n5022 VSS.n5020 204.757
R2231 VSS.n5022 VSS.n5021 204.757
R2232 VSS.n5029 VSS.n5028 204.757
R2233 VSS.n5030 VSS.n5029 204.757
R2234 VSS.n5030 VSS.n598 204.757
R2235 VSS.n5037 VSS.n598 204.757
R2236 VSS.n5038 VSS.n5037 204.757
R2237 VSS.n5039 VSS.n5038 204.757
R2238 VSS.n5042 VSS.n592 204.757
R2239 VSS.n5048 VSS.n592 204.757
R2240 VSS.n5049 VSS.n5048 204.757
R2241 VSS.n5051 VSS.n5049 204.757
R2242 VSS.n5051 VSS.n5050 204.757
R2243 VSS.n5058 VSS.n5057 204.757
R2244 VSS.n5060 VSS.n5058 204.757
R2245 VSS.n5060 VSS.n5059 204.757
R2246 VSS.n5059 VSS.n585 204.757
R2247 VSS.n5068 VSS.n585 204.757
R2248 VSS.n1190 VSS.n1189 200.845
R2249 VSS.n1051 VSS.n146 185
R2250 VSS.t85 VSS.n1051 185
R2251 VSS.n4168 VSS.n4167 185
R2252 VSS.n4170 VSS.n4169 185
R2253 VSS.n4172 VSS.n4171 185
R2254 VSS.n4174 VSS.n4173 185
R2255 VSS.n4176 VSS.n4175 185
R2256 VSS.n4178 VSS.n4177 185
R2257 VSS.n4179 VSS.n4160 185
R2258 VSS.t85 VSS.n4160 185
R2259 VSS.n4180 VSS.n4164 185
R2260 VSS.n5446 VSS.n5445 185
R2261 VSS.n5444 VSS.n5443 185
R2262 VSS.n5442 VSS.n142 185
R2263 VSS.n5440 VSS.n5439 185
R2264 VSS.n5438 VSS.n143 185
R2265 VSS.n5437 VSS.n5436 185
R2266 VSS.n5434 VSS.n144 185
R2267 VSS.n5432 VSS.n5431 185
R2268 VSS.n5430 VSS.n145 185
R2269 VSS.n145 VSS.t80 185
R2270 VSS.n3521 VSS.n101 185
R2271 VSS.t74 VSS.n101 185
R2272 VSS.n3520 VSS.n3519 185
R2273 VSS.n3518 VSS.n3517 185
R2274 VSS.n3516 VSS.n3515 185
R2275 VSS.n3514 VSS.n3513 185
R2276 VSS.n3512 VSS.n3511 185
R2277 VSS.n3510 VSS.n3509 185
R2278 VSS.n3508 VSS.n106 185
R2279 VSS.t74 VSS.n106 185
R2280 VSS.n3507 VSS.n110 185
R2281 VSS.n3608 VSS.n3607 185
R2282 VSS.n3604 VSS.n3603 185
R2283 VSS.n3602 VSS.n3601 185
R2284 VSS.n3600 VSS.n3599 185
R2285 VSS.n3598 VSS.n3597 185
R2286 VSS.n3596 VSS.n3595 185
R2287 VSS.n3594 VSS.n3593 185
R2288 VSS.n3592 VSS.n3591 185
R2289 VSS.n3548 VSS.n3522 185
R2290 VSS.t53 VSS.n3548 185
R2291 VSS.n3763 VSS.n3762 185
R2292 VSS.n3765 VSS.n3764 185
R2293 VSS.n3767 VSS.n3766 185
R2294 VSS.n3768 VSS.n3543 185
R2295 VSS.t53 VSS.n3543 185
R2296 VSS.n3770 VSS.n3769 185
R2297 VSS.n3772 VSS.n3771 185
R2298 VSS.n3774 VSS.n3773 185
R2299 VSS.n3776 VSS.n3775 185
R2300 VSS.n3777 VSS.n1114 185
R2301 VSS.n3625 VSS.n1216 185
R2302 VSS.n3627 VSS.n3626 185
R2303 VSS.n3628 VSS.n3620 185
R2304 VSS.n3630 VSS.n3629 185
R2305 VSS.n3632 VSS.n3618 185
R2306 VSS.n3634 VSS.n3633 185
R2307 VSS.n3635 VSS.n3617 185
R2308 VSS.n3637 VSS.n3636 185
R2309 VSS.n3637 VSS.t55 185
R2310 VSS.n3638 VSS.n3578 185
R2311 VSS.n3690 VSS.n1240 185
R2312 VSS.n3691 VSS.n3689 185
R2313 VSS.n3693 VSS.n3692 185
R2314 VSS.n3695 VSS.n3686 185
R2315 VSS.n3697 VSS.n3696 185
R2316 VSS.n3698 VSS.n3685 185
R2317 VSS.n3700 VSS.n3699 185
R2318 VSS.n3702 VSS.n3609 185
R2319 VSS.n3704 VSS.n3703 185
R2320 VSS.n3703 VSS.t55 185
R2321 VSS.n3430 VSS.n1274 185
R2322 VSS.n3432 VSS.n3431 185
R2323 VSS.n3433 VSS.n3428 185
R2324 VSS.n3435 VSS.n3434 185
R2325 VSS.n3437 VSS.n3427 185
R2326 VSS.n3438 VSS.n3426 185
R2327 VSS.n3441 VSS.n3440 185
R2328 VSS.n3442 VSS.n3424 185
R2329 VSS.n3424 VSS.t81 185
R2330 VSS.n3444 VSS.n3443 185
R2331 VSS.n3892 VSS.n3891 185
R2332 VSS.n3889 VSS.n1297 185
R2333 VSS.n3888 VSS.n3887 185
R2334 VSS.n3886 VSS.n3885 185
R2335 VSS.n3884 VSS.n1301 185
R2336 VSS.n3882 VSS.n3881 185
R2337 VSS.n3880 VSS.n1302 185
R2338 VSS.n3879 VSS.n3878 185
R2339 VSS.n3876 VSS.n1303 185
R2340 VSS.n3876 VSS.t81 185
R2341 VSS.n5075 VSS.n5074 185
R2342 VSS.n4693 VSS.n582 185
R2343 VSS.n4695 VSS.n4694 185
R2344 VSS.n4697 VSS.n4696 185
R2345 VSS.n4699 VSS.n4698 185
R2346 VSS.n4701 VSS.n4700 185
R2347 VSS.n4703 VSS.n4702 185
R2348 VSS.n4705 VSS.n4704 185
R2349 VSS.n4707 VSS.n4706 185
R2350 VSS.n733 VSS.n559 185
R2351 VSS.n732 VSS.n553 185
R2352 VSS.t73 VSS.n553 185
R2353 VSS.n731 VSS.n730 185
R2354 VSS.n729 VSS.n728 185
R2355 VSS.n727 VSS.n726 185
R2356 VSS.n725 VSS.n724 185
R2357 VSS.n723 VSS.n548 185
R2358 VSS.t73 VSS.n548 185
R2359 VSS.n722 VSS.n721 185
R2360 VSS.n668 VSS.n540 185
R2361 VSS.n4773 VSS.n4772 185
R2362 VSS.n4723 VSS.n4722 185
R2363 VSS.n4721 VSS.n4720 185
R2364 VSS.n4719 VSS.n4718 185
R2365 VSS.n4717 VSS.n4716 185
R2366 VSS.n4715 VSS.n4714 185
R2367 VSS.n4713 VSS.n4712 185
R2368 VSS.n4711 VSS.n4710 185
R2369 VSS.n4709 VSS.n4708 185
R2370 VSS.n4784 VSS.n536 185
R2371 VSS.n4785 VSS.n530 185
R2372 VSS.t76 VSS.n530 185
R2373 VSS.n4787 VSS.n4786 185
R2374 VSS.n4789 VSS.n4788 185
R2375 VSS.n4791 VSS.n4790 185
R2376 VSS.n4793 VSS.n4792 185
R2377 VSS.n4794 VSS.n525 185
R2378 VSS.t76 VSS.n525 185
R2379 VSS.n4796 VSS.n4795 185
R2380 VSS.n4799 VSS.n4798 185
R2381 VSS.n4806 VSS.n4803 185
R2382 VSS.n4808 VSS.n4807 185
R2383 VSS.n4809 VSS.n667 185
R2384 VSS.n4811 VSS.n4810 185
R2385 VSS.n4813 VSS.n666 185
R2386 VSS.n4814 VSS.n665 185
R2387 VSS.n4817 VSS.n4816 185
R2388 VSS.n4818 VSS.n663 185
R2389 VSS.n663 VSS.t79 185
R2390 VSS.n4820 VSS.n4819 185
R2391 VSS.n4883 VSS.n4882 185
R2392 VSS.n4885 VSS.n4836 185
R2393 VSS.n4887 VSS.n4886 185
R2394 VSS.n4888 VSS.n4835 185
R2395 VSS.n4890 VSS.n4889 185
R2396 VSS.n4892 VSS.n4833 185
R2397 VSS.n4894 VSS.n4893 185
R2398 VSS.n4895 VSS.n4830 185
R2399 VSS.n4897 VSS.n4896 185
R2400 VSS.n4897 VSS.t79 185
R2401 VSS.n1852 VSS.n1851 185
R2402 VSS.n1853 VSS.n1847 185
R2403 VSS.n1855 VSS.n1854 185
R2404 VSS.n1857 VSS.n1845 185
R2405 VSS.n1859 VSS.n1858 185
R2406 VSS.n1860 VSS.n1844 185
R2407 VSS.n1862 VSS.n1861 185
R2408 VSS.n1864 VSS.n1843 185
R2409 VSS.n1865 VSS.n1809 185
R2410 VSS.n1865 VSS.t75 185
R2411 VSS.n5160 VSS.n445 185
R2412 VSS.n5161 VSS.n444 185
R2413 VSS.n5164 VSS.n5163 185
R2414 VSS.n5165 VSS.n443 185
R2415 VSS.n443 VSS.t75 185
R2416 VSS.n5167 VSS.n5166 185
R2417 VSS.n5169 VSS.n441 185
R2418 VSS.n5171 VSS.n5170 185
R2419 VSS.n5172 VSS.n437 185
R2420 VSS.n5174 VSS.n5173 185
R2421 VSS.n831 VSS.n830 185
R2422 VSS.n829 VSS.n828 185
R2423 VSS.n827 VSS.n826 185
R2424 VSS.n825 VSS.n824 185
R2425 VSS.n823 VSS.n822 185
R2426 VSS.n821 VSS.n820 185
R2427 VSS.n819 VSS.n818 185
R2428 VSS.n817 VSS.n816 185
R2429 VSS.n815 VSS.n483 185
R2430 VSS.t58 VSS.n483 185
R2431 VSS.n4641 VSS.n744 185
R2432 VSS.n769 VSS.n745 185
R2433 VSS.n771 VSS.n770 185
R2434 VSS.n768 VSS.n757 185
R2435 VSS.n767 VSS.n766 185
R2436 VSS.n765 VSS.n764 185
R2437 VSS.n763 VSS.n762 185
R2438 VSS.n761 VSS.n760 185
R2439 VSS.n759 VSS.n758 185
R2440 VSS.n4602 VSS.n777 185
R2441 VSS.n4601 VSS.n773 185
R2442 VSS.t56 VSS.n773 185
R2443 VSS.n4600 VSS.n4599 185
R2444 VSS.n4598 VSS.n4597 185
R2445 VSS.n4596 VSS.n4595 185
R2446 VSS.n4594 VSS.n4593 185
R2447 VSS.n4592 VSS.n753 185
R2448 VSS.t56 VSS.n753 185
R2449 VSS.n4591 VSS.n4590 185
R2450 VSS.n4589 VSS.n4588 185
R2451 VSS.n3161 VSS.n3160 185
R2452 VSS.n3163 VSS.n3162 185
R2453 VSS.n3165 VSS.n3164 185
R2454 VSS.n3166 VSS.n478 185
R2455 VSS.t58 VSS.n478 185
R2456 VSS.n3168 VSS.n3167 185
R2457 VSS.n3170 VSS.n3169 185
R2458 VSS.n3172 VSS.n3171 185
R2459 VSS.n3174 VSS.n3173 185
R2460 VSS.n3176 VSS.n3175 185
R2461 VSS.n4506 VSS.n4505 185
R2462 VSS.n4462 VSS.n4461 185
R2463 VSS.n4460 VSS.n4459 185
R2464 VSS.n4458 VSS.n4457 185
R2465 VSS.n4456 VSS.n4455 185
R2466 VSS.n4454 VSS.n4453 185
R2467 VSS.n4452 VSS.n4451 185
R2468 VSS.n4450 VSS.n4449 185
R2469 VSS.n4448 VSS.n4447 185
R2470 VSS.n4423 VSS.n890 185
R2471 VSS.n4422 VSS.n884 185
R2472 VSS.t86 VSS.n884 185
R2473 VSS.n4421 VSS.n4420 185
R2474 VSS.n4419 VSS.n4418 185
R2475 VSS.n4417 VSS.n4416 185
R2476 VSS.n4415 VSS.n4414 185
R2477 VSS.n4413 VSS.n879 185
R2478 VSS.t86 VSS.n879 185
R2479 VSS.n4412 VSS.n4411 185
R2480 VSS.n4410 VSS.n869 185
R2481 VSS.n2397 VSS.n2396 185
R2482 VSS.n2376 VSS.n2375 185
R2483 VSS.n2374 VSS.n2063 185
R2484 VSS.n2372 VSS.n2371 185
R2485 VSS.n2370 VSS.n2064 185
R2486 VSS.n2369 VSS.n2368 185
R2487 VSS.n2366 VSS.n2065 185
R2488 VSS.n2364 VSS.n2363 185
R2489 VSS.n2362 VSS.n2066 185
R2490 VSS.n2066 VSS.t99 185
R2491 VSS.n4941 VSS.n638 185
R2492 VSS.n2377 VSS.n639 185
R2493 VSS.n2379 VSS.n2378 185
R2494 VSS.n2381 VSS.n2380 185
R2495 VSS.n2383 VSS.n2382 185
R2496 VSS.n2385 VSS.n2384 185
R2497 VSS.n2387 VSS.n2386 185
R2498 VSS.n2389 VSS.n2388 185
R2499 VSS.n2391 VSS.n2390 185
R2500 VSS.n2018 VSS.n656 185
R2501 VSS.n2019 VSS.n652 185
R2502 VSS.t96 VSS.n652 185
R2503 VSS.n2021 VSS.n2020 185
R2504 VSS.n2023 VSS.n2022 185
R2505 VSS.n2025 VSS.n2024 185
R2506 VSS.n2027 VSS.n2026 185
R2507 VSS.n2028 VSS.n647 185
R2508 VSS.t96 VSS.n647 185
R2509 VSS.n2030 VSS.n2029 185
R2510 VSS.n2032 VSS.n2031 185
R2511 VSS.n2433 VSS.n2017 185
R2512 VSS.n2435 VSS.n2434 185
R2513 VSS.n2437 VSS.n2016 185
R2514 VSS.n2438 VSS.n2015 185
R2515 VSS.n2438 VSS.t99 185
R2516 VSS.n2441 VSS.n2440 185
R2517 VSS.n2442 VSS.n2014 185
R2518 VSS.n2444 VSS.n2443 185
R2519 VSS.n2446 VSS.n2013 185
R2520 VSS.n2447 VSS.n2002 185
R2521 VSS.n2351 VSS.n2067 185
R2522 VSS.n2349 VSS.n2348 185
R2523 VSS.n2347 VSS.n2110 185
R2524 VSS.n2346 VSS.n2345 185
R2525 VSS.n2343 VSS.n2111 185
R2526 VSS.n2341 VSS.n2340 185
R2527 VSS.n2339 VSS.n2112 185
R2528 VSS.n2338 VSS.n2337 185
R2529 VSS.n2335 VSS.n2113 185
R2530 VSS.n2136 VSS.n2003 185
R2531 VSS.n2138 VSS.n2137 185
R2532 VSS.n2137 VSS.t71 185
R2533 VSS.n2140 VSS.n2139 185
R2534 VSS.n2142 VSS.n2134 185
R2535 VSS.n2144 VSS.n2143 185
R2536 VSS.n2146 VSS.n2145 185
R2537 VSS.n2147 VSS.n2132 185
R2538 VSS.n2147 VSS.t71 185
R2539 VSS.n2150 VSS.n2149 185
R2540 VSS.n2151 VSS.n2131 185
R2541 VSS.n2264 VSS.n1701 185
R2542 VSS.n2266 VSS.n2257 185
R2543 VSS.n2269 VSS.n2268 185
R2544 VSS.n2270 VSS.n2256 185
R2545 VSS.n2272 VSS.n2271 185
R2546 VSS.n2274 VSS.n2255 185
R2547 VSS.n2277 VSS.n2276 185
R2548 VSS.n2278 VSS.n2254 185
R2549 VSS.n2280 VSS.n2279 185
R2550 VSS.n2504 VSS.n2503 185
R2551 VSS.n2505 VSS.n1574 185
R2552 VSS.n1574 VSS.t98 185
R2553 VSS.n2507 VSS.n2506 185
R2554 VSS.n2509 VSS.n1573 185
R2555 VSS.n2511 VSS.n2510 185
R2556 VSS.n2513 VSS.n2512 185
R2557 VSS.n2514 VSS.n1571 185
R2558 VSS.n2514 VSS.t98 185
R2559 VSS.n2516 VSS.n2515 185
R2560 VSS.n2518 VSS.n2517 185
R2561 VSS.n3046 VSS.n1456 185
R2562 VSS.n1542 VSS.n1466 185
R2563 VSS.n1544 VSS.n1543 185
R2564 VSS.n1546 VSS.n1545 185
R2565 VSS.n1548 VSS.n1547 185
R2566 VSS.n1550 VSS.n1549 185
R2567 VSS.n1552 VSS.n1551 185
R2568 VSS.n1554 VSS.n1553 185
R2569 VSS.n1556 VSS.n1555 185
R2570 VSS.n2577 VSS.n1483 185
R2571 VSS.n2576 VSS.n1479 185
R2572 VSS.t84 VSS.n1479 185
R2573 VSS.n2575 VSS.n2574 185
R2574 VSS.n2573 VSS.n2572 185
R2575 VSS.n2571 VSS.n2570 185
R2576 VSS.n2569 VSS.n2568 185
R2577 VSS.n2567 VSS.n1474 185
R2578 VSS.t84 VSS.n1474 185
R2579 VSS.n2566 VSS.n2565 185
R2580 VSS.n2564 VSS.n2563 185
R2581 VSS.n5313 VSS.n328 185
R2582 VSS.n5311 VSS.n5310 185
R2583 VSS.n5309 VSS.n329 185
R2584 VSS.n5308 VSS.n5307 185
R2585 VSS.n5305 VSS.n330 185
R2586 VSS.n5303 VSS.n5302 185
R2587 VSS.n5301 VSS.n331 185
R2588 VSS.n5300 VSS.n5299 185
R2589 VSS.n5297 VSS.n332 185
R2590 VSS.n4371 VSS.n305 185
R2591 VSS.n4373 VSS.n4372 185
R2592 VSS.n4372 VSS.t78 185
R2593 VSS.n4375 VSS.n4374 185
R2594 VSS.n4377 VSS.n4370 185
R2595 VSS.n4379 VSS.n4378 185
R2596 VSS.n4381 VSS.n4380 185
R2597 VSS.n4382 VSS.n4368 185
R2598 VSS.n4382 VSS.t78 185
R2599 VSS.n4384 VSS.n4383 185
R2600 VSS.n4386 VSS.n4385 185
R2601 VSS.n4198 VSS.n4197 185
R2602 VSS.n4195 VSS.n4194 185
R2603 VSS.n4193 VSS.n4192 185
R2604 VSS.n4191 VSS.n4190 185
R2605 VSS.n4189 VSS.n4188 185
R2606 VSS.n4187 VSS.n4186 185
R2607 VSS.n4185 VSS.n4184 185
R2608 VSS.n4183 VSS.n4182 185
R2609 VSS.n4181 VSS.n1019 185
R2610 VSS.n2302 VSS.n2301 185
R2611 VSS.n2304 VSS.n2128 185
R2612 VSS.n2307 VSS.n2306 185
R2613 VSS.n2129 VSS.n2123 185
R2614 VSS.n2318 VSS.n2317 185
R2615 VSS.n2320 VSS.n2122 185
R2616 VSS.n2323 VSS.n2322 185
R2617 VSS.n2324 VSS.n2114 185
R2618 VSS.n2333 VSS.n2332 185
R2619 VSS.n2519 VSS.n1567 185
R2620 VSS.n2522 VSS.n2521 185
R2621 VSS.n2232 VSS.n1569 185
R2622 VSS.n2239 VSS.n2237 185
R2623 VSS.n2242 VSS.n2241 185
R2624 VSS.n2229 VSS.n2228 185
R2625 VSS.n2251 VSS.n2250 185
R2626 VSS.n2253 VSS.n2226 185
R2627 VSS.n2283 VSS.n2282 185
R2628 VSS.n2562 VSS.n2561 185
R2629 VSS.n1529 VSS.n1490 185
R2630 VSS.n1531 VSS.n1530 185
R2631 VSS.n2553 VSS.n2552 185
R2632 VSS.n2551 VSS.n2550 185
R2633 VSS.n1538 VSS.n1533 185
R2634 VSS.n1540 VSS.n1539 185
R2635 VSS.n2542 VSS.n2541 185
R2636 VSS.n2540 VSS.n2539 185
R2637 VSS.n4387 VSS.n4337 185
R2638 VSS.n4390 VSS.n4389 185
R2639 VSS.n4366 VSS.n4365 185
R2640 VSS.n4343 VSS.n4340 185
R2641 VSS.n4358 VSS.n4357 185
R2642 VSS.n4355 VSS.n4354 185
R2643 VSS.n4346 VSS.n4345 185
R2644 VSS.n4347 VSS.n333 185
R2645 VSS.n5295 VSS.n5294 185
R2646 VSS.n4103 VSS.n4102 185
R2647 VSS.n4075 VSS.n4068 185
R2648 VSS.n4077 VSS.n4076 185
R2649 VSS.n4094 VSS.n4093 185
R2650 VSS.n4092 VSS.n4091 185
R2651 VSS.n4081 VSS.n4079 185
R2652 VSS.n4083 VSS.n4082 185
R2653 VSS.n1018 VSS.n1016 185
R2654 VSS.n4322 VSS.n4321 185
R2655 VSS.n1981 VSS.n1980 185
R2656 VSS.n1983 VSS.n1982 185
R2657 VSS.n1985 VSS.n1984 185
R2658 VSS.n1987 VSS.n1986 185
R2659 VSS.n1989 VSS.n1988 185
R2660 VSS.n1991 VSS.n1990 185
R2661 VSS.n1993 VSS.n1992 185
R2662 VSS.n1995 VSS.n1994 185
R2663 VSS.n1996 VSS.n1607 185
R2664 VSS.t87 VSS.n1607 185
R2665 VSS.n1958 VSS.n1957 185
R2666 VSS.n1960 VSS.n1807 185
R2667 VSS.n1963 VSS.n1962 185
R2668 VSS.n1964 VSS.n1806 185
R2669 VSS.n1966 VSS.n1965 185
R2670 VSS.n1968 VSS.n1805 185
R2671 VSS.n1971 VSS.n1970 185
R2672 VSS.n1972 VSS.n1804 185
R2673 VSS.n1974 VSS.n1973 185
R2674 VSS.n1749 VSS.n1748 185
R2675 VSS.n1750 VSS.n1746 185
R2676 VSS.n1746 VSS.t83 185
R2677 VSS.n1752 VSS.n1751 185
R2678 VSS.n1754 VSS.n1745 185
R2679 VSS.n1756 VSS.n1755 185
R2680 VSS.n1758 VSS.n1757 185
R2681 VSS.n1759 VSS.n1743 185
R2682 VSS.n1759 VSS.t83 185
R2683 VSS.n1761 VSS.n1760 185
R2684 VSS.n1763 VSS.n1762 185
R2685 VSS.n1741 VSS.n1740 185
R2686 VSS.n1739 VSS.n1738 185
R2687 VSS.n1737 VSS.n1736 185
R2688 VSS.n1735 VSS.n1602 185
R2689 VSS.t87 VSS.n1602 185
R2690 VSS.n1734 VSS.n1733 185
R2691 VSS.n1732 VSS.n1731 185
R2692 VSS.n1730 VSS.n1729 185
R2693 VSS.n1728 VSS.n1727 185
R2694 VSS.n1726 VSS.n1725 185
R2695 VSS.n3073 VSS.n3072 185
R2696 VSS.n3071 VSS.n3070 185
R2697 VSS.n3069 VSS.n1452 185
R2698 VSS.n3067 VSS.n3066 185
R2699 VSS.n3065 VSS.n1453 185
R2700 VSS.n3064 VSS.n3063 185
R2701 VSS.n3061 VSS.n1454 185
R2702 VSS.n3059 VSS.n3058 185
R2703 VSS.n3057 VSS.n1455 185
R2704 VSS.n1455 VSS.t77 185
R2705 VSS.n3105 VSS.n1436 185
R2706 VSS.n3103 VSS.n3102 185
R2707 VSS.n3101 VSS.n1437 185
R2708 VSS.n3100 VSS.n3099 185
R2709 VSS.n3097 VSS.n1438 185
R2710 VSS.n3095 VSS.n3094 185
R2711 VSS.n3093 VSS.n1439 185
R2712 VSS.n3092 VSS.n3091 185
R2713 VSS.n3089 VSS.n1440 185
R2714 VSS.n2853 VSS.n2852 185
R2715 VSS.n2854 VSS.n2731 185
R2716 VSS.n2731 VSS.t68 185
R2717 VSS.n2856 VSS.n2855 185
R2718 VSS.n2858 VSS.n2730 185
R2719 VSS.n2860 VSS.n2859 185
R2720 VSS.n2862 VSS.n2861 185
R2721 VSS.n2863 VSS.n2728 185
R2722 VSS.n2863 VSS.t68 185
R2723 VSS.n2866 VSS.n2865 185
R2724 VSS.n2867 VSS.n2587 185
R2725 VSS.n2972 VSS.n2583 185
R2726 VSS.n2973 VSS.n2582 185
R2727 VSS.n2976 VSS.n2975 185
R2728 VSS.n2977 VSS.n2581 185
R2729 VSS.n2581 VSS.t77 185
R2730 VSS.n2979 VSS.n2978 185
R2731 VSS.n2981 VSS.n2579 185
R2732 VSS.n2983 VSS.n2982 185
R2733 VSS.n2984 VSS.n1487 185
R2734 VSS.n2986 VSS.n2985 185
R2735 VSS.n2717 VSS.n2622 185
R2736 VSS.n2715 VSS.n2714 185
R2737 VSS.n2713 VSS.n2673 185
R2738 VSS.n2712 VSS.n2711 185
R2739 VSS.n2709 VSS.n2674 185
R2740 VSS.n2707 VSS.n2706 185
R2741 VSS.n2705 VSS.n2675 185
R2742 VSS.n2704 VSS.n2703 185
R2743 VSS.n2701 VSS.n2676 185
R2744 VSS.n2701 VSS.t70 185
R2745 VSS.n239 VSS.n238 185
R2746 VSS.n2624 VSS.n2623 185
R2747 VSS.n2626 VSS.n2625 185
R2748 VSS.n2628 VSS.n2627 185
R2749 VSS.n2630 VSS.n2629 185
R2750 VSS.n2632 VSS.n2631 185
R2751 VSS.n2634 VSS.n2633 185
R2752 VSS.n2636 VSS.n2635 185
R2753 VSS.n2638 VSS.n2637 185
R2754 VSS.n3280 VSS.n189 185
R2755 VSS.n3279 VSS.n183 185
R2756 VSS.t59 VSS.n183 185
R2757 VSS.n3278 VSS.n3277 185
R2758 VSS.n3276 VSS.n3275 185
R2759 VSS.n3274 VSS.n3273 185
R2760 VSS.n3272 VSS.n3271 185
R2761 VSS.n3270 VSS.n178 185
R2762 VSS.t59 VSS.n178 185
R2763 VSS.n3269 VSS.n3268 185
R2764 VSS.n3267 VSS.n3266 185
R2765 VSS.n5331 VSS.n5330 185
R2766 VSS.n5333 VSS.n5332 185
R2767 VSS.n5335 VSS.n5328 185
R2768 VSS.n5336 VSS.n5327 185
R2769 VSS.n5336 VSS.t70 185
R2770 VSS.n5339 VSS.n5338 185
R2771 VSS.n5340 VSS.n5326 185
R2772 VSS.n5342 VSS.n5341 185
R2773 VSS.n5344 VSS.n5325 185
R2774 VSS.n5345 VSS.n306 185
R2775 VSS.n2719 VSS.n2718 185
R2776 VSS.n2671 VSS.n2670 185
R2777 VSS.n2648 VSS.n2647 185
R2778 VSS.n2662 VSS.n2661 185
R2779 VSS.n2659 VSS.n2658 185
R2780 VSS.n2650 VSS.n166 185
R2781 VSS.n5418 VSS.n5417 185
R2782 VSS.n5421 VSS.n5420 185
R2783 VSS.n165 VSS.n164 185
R2784 VSS.n3265 VSS.n161 185
R2785 VSS.n170 VSS.n162 185
R2786 VSS.n5416 VSS.n5415 185
R2787 VSS.n2651 VSS.n171 185
R2788 VSS.n2657 VSS.n2656 185
R2789 VSS.n2666 VSS.n2665 185
R2790 VSS.n2668 VSS.n2667 185
R2791 VSS.n2646 VSS.n2645 185
R2792 VSS.n2644 VSS.n2639 185
R2793 VSS.n3074 VSS.n1442 185
R2794 VSS.n3077 VSS.n3076 185
R2795 VSS.n2942 VSS.n1450 185
R2796 VSS.n2954 VSS.n2952 185
R2797 VSS.n2956 VSS.n2955 185
R2798 VSS.n2939 VSS.n2938 185
R2799 VSS.n2935 VSS.n2590 185
R2800 VSS.n2589 VSS.n2584 185
R2801 VSS.n2970 VSS.n2969 185
R2802 VSS.n2968 VSS.n2967 185
R2803 VSS.n2965 VSS.n2964 185
R2804 VSS.n2936 VSS.n2588 185
R2805 VSS.n2947 VSS.n2932 185
R2806 VSS.n2948 VSS.n2933 185
R2807 VSS.n2951 VSS.n2950 185
R2808 VSS.n2945 VSS.n1447 185
R2809 VSS.n1449 VSS.n1441 185
R2810 VSS.n3087 VSS.n3086 185
R2811 VSS.n1979 VSS.n1978 185
R2812 VSS.n1711 VSS.n1710 185
R2813 VSS.n1709 VSS.n1708 185
R2814 VSS.n1790 VSS.n1789 185
R2815 VSS.n1788 VSS.n1787 185
R2816 VSS.n1777 VSS.n1776 185
R2817 VSS.n1775 VSS.n1774 185
R2818 VSS.n1770 VSS.n1769 185
R2819 VSS.n1768 VSS.n1767 185
R2820 VSS.n1766 VSS.n1765 185
R2821 VSS.n1771 VSS.n1719 185
R2822 VSS.n1781 VSS.n1780 185
R2823 VSS.n1783 VSS.n1718 185
R2824 VSS.n1786 VSS.n1785 185
R2825 VSS.n1791 VSS.n1707 185
R2826 VSS.n1801 VSS.n1800 185
R2827 VSS.n1803 VSS.n1706 185
R2828 VSS.n1977 VSS.n1976 185
R2829 VSS.n2399 VSS.n2398 185
R2830 VSS.n2056 VSS.n2050 185
R2831 VSS.n2410 VSS.n2409 185
R2832 VSS.n2412 VSS.n2049 185
R2833 VSS.n2414 VSS.n2413 185
R2834 VSS.n2043 VSS.n2037 185
R2835 VSS.n2425 VSS.n2424 185
R2836 VSS.n2427 VSS.n2036 185
R2837 VSS.n2429 VSS.n2428 185
R2838 VSS.n2034 VSS.n2033 185
R2839 VSS.n2421 VSS.n2420 185
R2840 VSS.n2423 VSS.n2422 185
R2841 VSS.n2045 VSS.n2044 185
R2842 VSS.n2047 VSS.n2046 185
R2843 VSS.n2406 VSS.n2405 185
R2844 VSS.n2408 VSS.n2407 185
R2845 VSS.n2058 VSS.n2057 185
R2846 VSS.n2060 VSS.n2059 185
R2847 VSS.n3140 VSS.n1389 185
R2848 VSS.n3138 VSS.n3137 185
R2849 VSS.n3136 VSS.n1417 185
R2850 VSS.n3135 VSS.n3134 185
R2851 VSS.n3132 VSS.n1418 185
R2852 VSS.n3130 VSS.n3129 185
R2853 VSS.n3128 VSS.n1419 185
R2854 VSS.n3127 VSS.n3126 185
R2855 VSS.n3124 VSS.n1420 185
R2856 VSS.n3124 VSS.t100 185
R2857 VSS.n4541 VSS.n847 185
R2858 VSS.n1390 VSS.n848 185
R2859 VSS.n1392 VSS.n1391 185
R2860 VSS.n1394 VSS.n1393 185
R2861 VSS.n1396 VSS.n1395 185
R2862 VSS.n1398 VSS.n1397 185
R2863 VSS.n1400 VSS.n1399 185
R2864 VSS.n1402 VSS.n1401 185
R2865 VSS.n1404 VSS.n1403 185
R2866 VSS.n899 VSS.n865 185
R2867 VSS.n2775 VSS.n861 185
R2868 VSS.t88 VSS.n861 185
R2869 VSS.n2777 VSS.n2776 185
R2870 VSS.n2779 VSS.n2778 185
R2871 VSS.n2781 VSS.n2780 185
R2872 VSS.n2783 VSS.n2782 185
R2873 VSS.n2784 VSS.n856 185
R2874 VSS.t88 VSS.n856 185
R2875 VSS.n2786 VSS.n2785 185
R2876 VSS.n2788 VSS.n2787 185
R2877 VSS.n2794 VSS.n2742 185
R2878 VSS.n2795 VSS.n2741 185
R2879 VSS.n2798 VSS.n2797 185
R2880 VSS.n2799 VSS.n2740 185
R2881 VSS.n2740 VSS.t100 185
R2882 VSS.n2801 VSS.n2800 185
R2883 VSS.n2803 VSS.n2738 185
R2884 VSS.n2805 VSS.n2804 185
R2885 VSS.n2806 VSS.n2737 185
R2886 VSS.n2808 VSS.n2807 185
R2887 VSS.n1341 VSS.n1340 185
R2888 VSS.n1338 VSS.n1337 185
R2889 VSS.n1336 VSS.n1335 185
R2890 VSS.n1334 VSS.n1333 185
R2891 VSS.n1332 VSS.n1331 185
R2892 VSS.n1330 VSS.n1329 185
R2893 VSS.n1328 VSS.n1327 185
R2894 VSS.n1326 VSS.n1325 185
R2895 VSS.n240 VSS.n217 185
R2896 VSS.t95 VSS.n217 185
R2897 VSS.n3859 VSS.n1318 185
R2898 VSS.n3857 VSS.n3856 185
R2899 VSS.n3855 VSS.n1319 185
R2900 VSS.n3854 VSS.n3853 185
R2901 VSS.n3851 VSS.n1320 185
R2902 VSS.n3849 VSS.n3848 185
R2903 VSS.n3847 VSS.n1321 185
R2904 VSS.n3846 VSS.n3845 185
R2905 VSS.n3843 VSS.n1322 185
R2906 VSS.n3481 VSS.n3418 185
R2907 VSS.n3482 VSS.n3417 185
R2908 VSS.n3482 VSS.t82 185
R2909 VSS.n3484 VSS.n3483 185
R2910 VSS.n3486 VSS.n3485 185
R2911 VSS.n3487 VSS.n3415 185
R2912 VSS.n3490 VSS.n3489 185
R2913 VSS.n3491 VSS.n3414 185
R2914 VSS.n3414 VSS.t82 185
R2915 VSS.n3493 VSS.n3492 185
R2916 VSS.n3495 VSS.n3264 185
R2917 VSS.n3366 VSS.n3365 185
R2918 VSS.n3364 VSS.n3363 185
R2919 VSS.n3362 VSS.n3361 185
R2920 VSS.n3360 VSS.n212 185
R2921 VSS.t95 VSS.n212 185
R2922 VSS.n3359 VSS.n3358 185
R2923 VSS.n3357 VSS.n3356 185
R2924 VSS.n3355 VSS.n3354 185
R2925 VSS.n3353 VSS.n3352 185
R2926 VSS.n3351 VSS.n3350 185
R2927 VSS.n1339 VSS.n1324 185
R2928 VSS.n3389 VSS.n3388 185
R2929 VSS.n3387 VSS.n3386 185
R2930 VSS.n3404 VSS.n3403 185
R2931 VSS.n3406 VSS.n3405 185
R2932 VSS.n3377 VSS.n3376 185
R2933 VSS.n3375 VSS.n3374 185
R2934 VSS.n3501 VSS.n3500 185
R2935 VSS.n3503 VSS.n3502 185
R2936 VSS.n3496 VSS.n3367 185
R2937 VSS.n3499 VSS.n3498 185
R2938 VSS.n3413 VSS.n3412 185
R2939 VSS.n3398 VSS.n3378 185
R2940 VSS.n3399 VSS.n3379 185
R2941 VSS.n3402 VSS.n3401 185
R2942 VSS.n3397 VSS.n3396 185
R2943 VSS.n3390 VSS.n1323 185
R2944 VSS.n3841 VSS.n3840 185
R2945 VSS.n3141 VSS.n1405 185
R2946 VSS.n3143 VSS.n1406 185
R2947 VSS.n3145 VSS.n3144 185
R2948 VSS.n2755 VSS.n2752 185
R2949 VSS.n2761 VSS.n2760 185
R2950 VSS.n2764 VSS.n2763 185
R2951 VSS.n2751 VSS.n2748 185
R2952 VSS.n2771 VSS.n2743 185
R2953 VSS.n2792 VSS.n2791 185
R2954 VSS.n2790 VSS.n2789 185
R2955 VSS.n2770 VSS.n2769 185
R2956 VSS.n2768 VSS.n2767 185
R2957 VSS.n2757 VSS.n2749 185
R2958 VSS.n2759 VSS.n2758 185
R2959 VSS.n1413 VSS.n1411 185
R2960 VSS.n1415 VSS.n1414 185
R2961 VSS.n3154 VSS.n3153 185
R2962 VSS.n3156 VSS.n3155 185
R2963 VSS.n4543 VSS.n4542 185
R2964 VSS.n924 VSS.n923 185
R2965 VSS.n926 VSS.n925 185
R2966 VSS.n917 VSS.n916 185
R2967 VSS.n915 VSS.n911 185
R2968 VSS.n938 VSS.n937 185
R2969 VSS.n940 VSS.n939 185
R2970 VSS.n905 VSS.n866 185
R2971 VSS.n4538 VSS.n4537 185
R2972 VSS.n4536 VSS.n4535 185
R2973 VSS.n906 VSS.n870 185
R2974 VSS.n908 VSS.n907 185
R2975 VSS.n936 VSS.n935 185
R2976 VSS.n934 VSS.n933 185
R2977 VSS.n919 VSS.n918 185
R2978 VSS.n921 VSS.n920 185
R2979 VSS.n873 VSS.n844 185
R2980 VSS.n872 VSS.n845 185
R2981 VSS.n833 VSS.n832 185
R2982 VSS.n4565 VSS.n4564 185
R2983 VSS.n4567 VSS.n4566 185
R2984 VSS.n808 VSS.n807 185
R2985 VSS.n806 VSS.n800 185
R2986 VSS.n4578 VSS.n4577 185
R2987 VSS.n4580 VSS.n4579 185
R2988 VSS.n790 VSS.n789 185
R2989 VSS.n788 VSS.n787 185
R2990 VSS.n4587 VSS.n4586 185
R2991 VSS.n795 VSS.n794 185
R2992 VSS.n797 VSS.n796 185
R2993 VSS.n4576 VSS.n4575 185
R2994 VSS.n4574 VSS.n4573 185
R2995 VSS.n810 VSS.n809 185
R2996 VSS.n812 VSS.n811 185
R2997 VSS.n4563 VSS.n4562 185
R2998 VSS.n4561 VSS.n4560 185
R2999 VSS.n1850 VSS.n484 185
R3000 VSS.n493 VSS.n466 185
R3001 VSS.n5141 VSS.n5140 185
R3002 VSS.n5143 VSS.n465 185
R3003 VSS.n5145 VSS.n5144 185
R3004 VSS.n463 VSS.n462 185
R3005 VSS.n461 VSS.n452 185
R3006 VSS.n451 VSS.n446 185
R3007 VSS.n5158 VSS.n5157 185
R3008 VSS.n5156 VSS.n5155 185
R3009 VSS.n5154 VSS.n5153 185
R3010 VSS.n5131 VSS.n5130 185
R3011 VSS.n5132 VSS.n458 185
R3012 VSS.n5134 VSS.n459 185
R3013 VSS.n5136 VSS.n5135 185
R3014 VSS.n5139 VSS.n5138 185
R3015 VSS.n494 VSS.n469 185
R3016 VSS.n5128 VSS.n5127 185
R3017 VSS.n4839 VSS.n4838 185
R3018 VSS.n4854 VSS.n4840 185
R3019 VSS.n4855 VSS.n4841 185
R3020 VSS.n4858 VSS.n4857 185
R3021 VSS.n4852 VSS.n4851 185
R3022 VSS.n4845 VSS.n513 185
R3023 VSS.n5113 VSS.n5112 185
R3024 VSS.n5116 VSS.n5115 185
R3025 VSS.n4800 VSS.n512 185
R3026 VSS.n4797 VSS.n510 185
R3027 VSS.n517 VSS.n511 185
R3028 VSS.n5111 VSS.n5110 185
R3029 VSS.n4846 VSS.n518 185
R3030 VSS.n4843 VSS.n4842 185
R3031 VSS.n4865 VSS.n4864 185
R3032 VSS.n4867 VSS.n4866 185
R3033 VSS.n4874 VSS.n4873 185
R3034 VSS.n4876 VSS.n4875 185
R3035 VSS.n4771 VSS.n4770 185
R3036 VSS.n4765 VSS.n4764 185
R3037 VSS.n4763 VSS.n4762 185
R3038 VSS.n4757 VSS.n4756 185
R3039 VSS.n4755 VSS.n4754 185
R3040 VSS.n4749 VSS.n4748 185
R3041 VSS.n4747 VSS.n4746 185
R3042 VSS.n4729 VSS.n537 185
R3043 VSS.n5107 VSS.n5106 185
R3044 VSS.n5105 VSS.n5104 185
R3045 VSS.n4730 VSS.n541 185
R3046 VSS.n4745 VSS.n4744 185
R3047 VSS.n4751 VSS.n4750 185
R3048 VSS.n4753 VSS.n4752 185
R3049 VSS.n4759 VSS.n4758 185
R3050 VSS.n4761 VSS.n4760 185
R3051 VSS.n4768 VSS.n4767 185
R3052 VSS.n4766 VSS.n4692 185
R3053 VSS.n5077 VSS.n5076 185
R3054 VSS.n580 VSS.n579 185
R3055 VSS.n578 VSS.n571 185
R3056 VSS.n5086 VSS.n5085 185
R3057 VSS.n5088 VSS.n5087 185
R3058 VSS.n5092 VSS.n5091 185
R3059 VSS.n5090 VSS.n569 185
R3060 VSS.n562 VSS.n560 185
R3061 VSS.n5101 VSS.n5100 185
R3062 VSS.n4643 VSS.n4642 185
R3063 VSS.n4614 VSS.n740 185
R3064 VSS.n4616 VSS.n4615 185
R3065 VSS.n4623 VSS.n4622 185
R3066 VSS.n4625 VSS.n4624 185
R3067 VSS.n4629 VSS.n4628 185
R3068 VSS.n4627 VSS.n4611 185
R3069 VSS.n780 VSS.n778 185
R3070 VSS.n4638 VSS.n4637 185
R3071 VSS.n4508 VSS.n4507 185
R3072 VSS.n4443 VSS.n4442 185
R3073 VSS.n4441 VSS.n4434 185
R3074 VSS.n4517 VSS.n4516 185
R3075 VSS.n4519 VSS.n4518 185
R3076 VSS.n4523 VSS.n4522 185
R3077 VSS.n4521 VSS.n4432 185
R3078 VSS.n893 VSS.n891 185
R3079 VSS.n4532 VSS.n4531 185
R3080 VSS.n1299 VSS.n1296 185
R3081 VSS.n1288 VSS.n1286 185
R3082 VSS.n3934 VSS.n3933 185
R3083 VSS.n3936 VSS.n1285 185
R3084 VSS.n3938 VSS.n3937 185
R3085 VSS.n1280 VSS.n1278 185
R3086 VSS.n3949 VSS.n3948 185
R3087 VSS.n3951 VSS.n1277 185
R3088 VSS.n3953 VSS.n3952 185
R3089 VSS.n3967 VSS.n3966 185
R3090 VSS.n3970 VSS.n3969 185
R3091 VSS.n1239 VSS.n1236 185
R3092 VSS.n1234 VSS.n1227 185
R3093 VSS.n3979 VSS.n3978 185
R3094 VSS.n3981 VSS.n1226 185
R3095 VSS.n3983 VSS.n3982 185
R3096 VSS.n3622 VSS.n1223 185
R3097 VSS.n3623 VSS.n1217 185
R3098 VSS.n3606 VSS.n3605 185
R3099 VSS.n3680 VSS.n3679 185
R3100 VSS.n3678 VSS.n3677 185
R3101 VSS.n3670 VSS.n3669 185
R3102 VSS.n3668 VSS.n3667 185
R3103 VSS.n3661 VSS.n3660 185
R3104 VSS.n3659 VSS.n3658 185
R3105 VSS.n3652 VSS.n3651 185
R3106 VSS.n3650 VSS.n3580 185
R3107 VSS.n3649 VSS.n3648 185
R3108 VSS.n3647 VSS.n3616 185
R3109 VSS.n3645 VSS.n3615 185
R3110 VSS.n3644 VSS.n3614 185
R3111 VSS.n3642 VSS.n3613 185
R3112 VSS.n3641 VSS.n3612 185
R3113 VSS.n3676 VSS.n3610 185
R3114 VSS.n3682 VSS.n3681 185
R3115 VSS.n3684 VSS.n3590 185
R3116 VSS.n3860 VSS.n1309 185
R3117 VSS.n3862 VSS.n1308 185
R3118 VSS.n3864 VSS.n3863 185
R3119 VSS.n3456 VSS.n3453 185
R3120 VSS.n3467 VSS.n3466 185
R3121 VSS.n3469 VSS.n3452 185
R3122 VSS.n3471 VSS.n3470 185
R3123 VSS.n3447 VSS.n3419 185
R3124 VSS.n3479 VSS.n3478 185
R3125 VSS.n3477 VSS.n3476 185
R3126 VSS.n3475 VSS.n3474 185
R3127 VSS.n3460 VSS.n3448 185
R3128 VSS.n3462 VSS.n3461 185
R3129 VSS.n3465 VSS.n3464 185
R3130 VSS.n3459 VSS.n1314 185
R3131 VSS.n1316 VSS.n1307 185
R3132 VSS.n3873 VSS.n3872 185
R3133 VSS.n3875 VSS.n1306 185
R3134 VSS.n3563 VSS.n3562 185
R3135 VSS.n3569 VSS.n3568 185
R3136 VSS.n3571 VSS.n3570 185
R3137 VSS.n3558 VSS.n3557 185
R3138 VSS.n3556 VSS.n3555 185
R3139 VSS.n3790 VSS.n3789 185
R3140 VSS.n3792 VSS.n3791 185
R3141 VSS.n3781 VSS.n3780 185
R3142 VSS.n3779 VSS.n1116 185
R3143 VSS.n3784 VSS.n3783 185
R3144 VSS.n3778 VSS.n3527 185
R3145 VSS.n3533 VSS.n3528 185
R3146 VSS.n3788 VSS.n3787 185
R3147 VSS.n3554 VSS.n3534 185
R3148 VSS.n3575 VSS.n3574 185
R3149 VSS.n3559 VSS.n3551 185
R3150 VSS.n3567 VSS.n3566 185
R3151 VSS.n3549 VSS.n3523 185
R3152 VSS.n4026 VSS.n4025 185
R3153 VSS.n4028 VSS.n4027 185
R3154 VSS.n4030 VSS.n4029 185
R3155 VSS.n4032 VSS.n4031 185
R3156 VSS.n4034 VSS.n4033 185
R3157 VSS.n4036 VSS.n4035 185
R3158 VSS.n4038 VSS.n4037 185
R3159 VSS.n4040 VSS.n4039 185
R3160 VSS.n4043 VSS.n4042 185
R3161 VSS.n4047 VSS.n1113 185
R3162 VSS.n4049 VSS.n4048 185
R3163 VSS.n4051 VSS.n1111 185
R3164 VSS.n4052 VSS.n1110 185
R3165 VSS.n4052 VSS.t80 185
R3166 VSS.n4055 VSS.n4054 185
R3167 VSS.n4056 VSS.n1109 185
R3168 VSS.n4058 VSS.n4057 185
R3169 VSS.n4060 VSS.n1108 185
R3170 VSS.n4063 VSS.n4062 185
R3171 VSS.n4943 VSS.n4942 185
R3172 VSS.n4906 VSS.n4905 185
R3173 VSS.n4908 VSS.n4907 185
R3174 VSS.n4915 VSS.n4914 185
R3175 VSS.n4913 VSS.n4829 185
R3176 VSS.n4927 VSS.n4926 185
R3177 VSS.n4925 VSS.n4824 185
R3178 VSS.n4823 VSS.n657 185
R3179 VSS.n4938 VSS.n4937 185
R3180 VSS.n4936 VSS.n4935 185
R3181 VSS.n4934 VSS.n4933 185
R3182 VSS.n4827 VSS.n4825 185
R3183 VSS.n4924 VSS.n4923 185
R3184 VSS.n4921 VSS.n4920 185
R3185 VSS.n4912 VSS.n4828 185
R3186 VSS.n4903 VSS.n4902 185
R3187 VSS.n4900 VSS.n635 185
R3188 VSS.n4898 VSS.n636 185
R3189 VSS.n1870 VSS.n1808 185
R3190 VSS.n1834 VSS.n1815 185
R3191 VSS.n1836 VSS.n1835 185
R3192 VSS.n1831 VSS.n1830 185
R3193 VSS.n1826 VSS.n1821 185
R3194 VSS.n1822 VSS.n432 185
R3195 VSS.n5182 VSS.n5181 185
R3196 VSS.n5185 VSS.n5184 185
R3197 VSS.n438 VSS.n431 185
R3198 VSS.n5176 VSS.n429 185
R3199 VSS.n5177 VSS.n430 185
R3200 VSS.n5180 VSS.n5179 185
R3201 VSS.n1823 VSS.n436 185
R3202 VSS.n1827 VSS.n1819 185
R3203 VSS.n1840 VSS.n1839 185
R3204 VSS.n1842 VSS.n1817 185
R3205 VSS.n1869 VSS.n1868 185
R3206 VSS.n1866 VSS.n1810 185
R3207 VSS.n3106 VSS.n1424 185
R3208 VSS.n3108 VSS.n1423 185
R3209 VSS.n3110 VSS.n3109 185
R3210 VSS.n2835 VSS.n2834 185
R3211 VSS.n2837 VSS.n2836 185
R3212 VSS.n2831 VSS.n2830 185
R3213 VSS.n2821 VSS.n2812 185
R3214 VSS.n2811 VSS.n2734 185
R3215 VSS.n2850 VSS.n2849 185
R3216 VSS.n2848 VSS.n2847 185
R3217 VSS.n2846 VSS.n2845 185
R3218 VSS.n2828 VSS.n2827 185
R3219 VSS.n2826 VSS.n2818 185
R3220 VSS.n2824 VSS.n2819 185
R3221 VSS.n2823 VSS.n1429 185
R3222 VSS.n1431 VSS.n1422 185
R3223 VSS.n3121 VSS.n3120 185
R3224 VSS.n3123 VSS.n1421 185
R3225 VSS.n237 VSS.n233 185
R3226 VSS.n5387 VSS.n5386 185
R3227 VSS.n5385 VSS.n220 185
R3228 VSS.n227 VSS.n226 185
R3229 VSS.n225 VSS.n224 185
R3230 VSS.n5401 VSS.n5400 185
R3231 VSS.n5399 VSS.n196 185
R3232 VSS.n195 VSS.n190 185
R3233 VSS.n5412 VSS.n5411 185
R3234 VSS.n5410 VSS.n5409 185
R3235 VSS.n5408 VSS.n5407 185
R3236 VSS.n202 VSS.n200 185
R3237 VSS.n5398 VSS.n5397 185
R3238 VSS.n223 VSS.n203 185
R3239 VSS.n5394 VSS.n5393 185
R3240 VSS.n232 VSS.n219 185
R3241 VSS.n5384 VSS.n5383 185
R3242 VSS.n236 VSS.n235 185
R3243 VSS.n5447 VSS.n112 185
R3244 VSS.n5450 VSS.n5449 185
R3245 VSS.n140 VSS.n139 185
R3246 VSS.n134 VSS.n133 185
R3247 VSS.n132 VSS.n131 185
R3248 VSS.n123 VSS.n87 185
R3249 VSS.n5466 VSS.n5465 185
R3250 VSS.n5469 VSS.n5468 185
R3251 VSS.n4044 VSS.n86 185
R3252 VSS.n4041 VSS.n84 185
R3253 VSS.n91 VSS.n85 185
R3254 VSS.n5464 VSS.n5463 185
R3255 VSS.n124 VSS.n92 185
R3256 VSS.n130 VSS.n129 185
R3257 VSS.n136 VSS.n135 185
R3258 VSS.n138 VSS.n137 185
R3259 VSS.n5451 VSS.n111 185
R3260 VSS.n5460 VSS.n5459 185
R3261 VSS.n1102 VSS.n1101 185
R3262 VSS.n1075 VSS.n1074 185
R3263 VSS.n1077 VSS.n1076 185
R3264 VSS.n1087 VSS.n1086 185
R3265 VSS.n1085 VSS.n1084 185
R3266 VSS.n1079 VSS.n1056 185
R3267 VSS.n4158 VSS.n4157 185
R3268 VSS.n4151 VSS.n1055 185
R3269 VSS.n4140 VSS.n4139 185
R3270 VSS.n1061 VSS.n1060 185
R3271 VSS.n4153 VSS.n4152 185
R3272 VSS.n4156 VSS.n4155 185
R3273 VSS.n1080 VSS.n1059 185
R3274 VSS.n1078 VSS.n1071 185
R3275 VSS.n1094 VSS.n1093 185
R3276 VSS.n1096 VSS.n1069 185
R3277 VSS.n1097 VSS.n1068 185
R3278 VSS.n1100 VSS.n1099 185
R3279 VSS.n4137 VSS.n4136 185
R3280 VSS.n4135 VSS.n4134 185
R3281 VSS.n4133 VSS.n4132 185
R3282 VSS.n4131 VSS.n4130 185
R3283 VSS.n4129 VSS.n4128 185
R3284 VSS.n4127 VSS.n4126 185
R3285 VSS.n4125 VSS.n4124 185
R3286 VSS.n4123 VSS.n4122 185
R3287 VSS.n4121 VSS.n1041 185
R3288 VSS.n4118 VSS.n1037 185
R3289 VSS.n4117 VSS.n1031 185
R3290 VSS.t97 VSS.n1031 185
R3291 VSS.n4116 VSS.n4115 185
R3292 VSS.n4114 VSS.n4113 185
R3293 VSS.n4112 VSS.n4111 185
R3294 VSS.n4110 VSS.n4109 185
R3295 VSS.n4108 VSS.n1026 185
R3296 VSS.t97 VSS.n1026 185
R3297 VSS.n4107 VSS.n4106 185
R3298 VSS.n4105 VSS.n4104 185
R3299 VSS.n2353 VSS.n2352 185
R3300 VSS.n2108 VSS.n2107 185
R3301 VSS.n2078 VSS.n2077 185
R3302 VSS.n2097 VSS.n2096 185
R3303 VSS.n2094 VSS.n2093 185
R3304 VSS.n2085 VSS.n2009 185
R3305 VSS.n2455 VSS.n2454 185
R3306 VSS.n2458 VSS.n2457 185
R3307 VSS.n2008 VSS.n2004 185
R3308 VSS.n2449 VSS.n2006 185
R3309 VSS.n2450 VSS.n2007 185
R3310 VSS.n2453 VSS.n2452 185
R3311 VSS.n2086 VSS.n2012 185
R3312 VSS.n2092 VSS.n2083 185
R3313 VSS.n2102 VSS.n2101 185
R3314 VSS.n2105 VSS.n2104 185
R3315 VSS.n2081 VSS.n2076 185
R3316 VSS.n2079 VSS.n2068 185
R3317 VSS.n2263 VSS.n2262 185
R3318 VSS.n2260 VSS.n1611 185
R3319 VSS.n2259 VSS.n1610 185
R3320 VSS.n1690 VSS.n1590 185
R3321 VSS.n2487 VSS.n2486 185
R3322 VSS.n2490 VSS.n2489 185
R3323 VSS.n1589 VSS.n1582 185
R3324 VSS.n1581 VSS.n1576 185
R3325 VSS.n2501 VSS.n2500 185
R3326 VSS.n2499 VSS.n2498 185
R3327 VSS.n2497 VSS.n2496 185
R3328 VSS.n2481 VSS.n1586 185
R3329 VSS.n2482 VSS.n1587 185
R3330 VSS.n2485 VSS.n2484 185
R3331 VSS.n1691 VSS.n1593 185
R3332 VSS.n2479 VSS.n2478 185
R3333 VSS.n1696 VSS.n1609 185
R3334 VSS.n1700 VSS.n1699 185
R3335 VSS.n3048 VSS.n3047 185
R3336 VSS.n3020 VSS.n3019 185
R3337 VSS.n3018 VSS.n3017 185
R3338 VSS.n3028 VSS.n3027 185
R3339 VSS.n3030 VSS.n3029 185
R3340 VSS.n3007 VSS.n3006 185
R3341 VSS.n3005 VSS.n2990 185
R3342 VSS.n2989 VSS.n1484 185
R3343 VSS.n3043 VSS.n3042 185
R3344 VSS.n3041 VSS.n3040 185
R3345 VSS.n3039 VSS.n3038 185
R3346 VSS.n3010 VSS.n3009 185
R3347 VSS.n3011 VSS.n2998 185
R3348 VSS.n3013 VSS.n2999 185
R3349 VSS.n3026 VSS.n3025 185
R3350 VSS.n3023 VSS.n3022 185
R3351 VSS.n3016 VSS.n1463 185
R3352 VSS.n3014 VSS.n1464 185
R3353 VSS.n5315 VSS.n5314 185
R3354 VSS.n2689 VSS.n2688 185
R3355 VSS.n2691 VSS.n2690 185
R3356 VSS.n2685 VSS.n2684 185
R3357 VSS.n2680 VSS.n315 185
R3358 VSS.n314 VSS.n310 185
R3359 VSS.n5354 VSS.n5353 185
R3360 VSS.n5356 VSS.n309 185
R3361 VSS.n5358 VSS.n5357 185
R3362 VSS.n5347 VSS.n307 185
R3363 VSS.n5349 VSS.n5348 185
R3364 VSS.n5352 VSS.n5351 185
R3365 VSS.n5324 VSS.n5323 185
R3366 VSS.n2681 VSS.n2678 185
R3367 VSS.n2695 VSS.n2694 185
R3368 VSS.n2697 VSS.n2677 185
R3369 VSS.n2698 VSS.n323 185
R3370 VSS.n2700 VSS.n326 185
R3371 VSS.n4196 VSS.n4166 185
R3372 VSS.n4302 VSS.n4301 185
R3373 VSS.n4300 VSS.n4299 185
R3374 VSS.n4294 VSS.n4293 185
R3375 VSS.n4292 VSS.n4291 185
R3376 VSS.n4286 VSS.n4285 185
R3377 VSS.n4284 VSS.n4283 185
R3378 VSS.n4266 VSS.n1038 185
R3379 VSS.n4318 VSS.n4317 185
R3380 VSS.n4316 VSS.n4315 185
R3381 VSS.n4267 VSS.n1042 185
R3382 VSS.n4282 VSS.n4281 185
R3383 VSS.n4288 VSS.n4287 185
R3384 VSS.n4290 VSS.n4289 185
R3385 VSS.n4296 VSS.n4295 185
R3386 VSS.n4298 VSS.n4297 185
R3387 VSS.n4303 VSS.n4165 185
R3388 VSS.n4312 VSS.n4311 185
R3389 VSS.n5564 VSS.n4 180.513
R3390 VSS.n5566 VSS.n5565 176.267
R3391 VSS.n4069 VSS.n6 175.546
R3392 VSS.n4100 VSS.n4069 175.546
R3393 VSS.n4100 VSS.n4070 175.546
R3394 VSS.n4096 VSS.n4070 175.546
R3395 VSS.n4096 VSS.n4073 175.546
R3396 VSS.n4089 VSS.n4073 175.546
R3397 VSS.n4089 VSS.n4085 175.546
R3398 VSS.n4085 VSS.n1015 175.546
R3399 VSS.n4324 VSS.n1015 175.546
R3400 VSS.n4324 VSS.n1014 175.546
R3401 VSS.n4328 VSS.n1014 175.546
R3402 VSS.n5560 VSS.n5559 175.546
R3403 VSS.n5559 VSS.n8 175.546
R3404 VSS.n5555 VSS.n8 175.546
R3405 VSS.n5555 VSS.n10 175.546
R3406 VSS.n5551 VSS.n10 175.546
R3407 VSS.n5551 VSS.n13 175.546
R3408 VSS.n5547 VSS.n13 175.546
R3409 VSS.n5547 VSS.n27 175.546
R3410 VSS.n5543 VSS.n27 175.546
R3411 VSS.n5543 VSS.n29 175.546
R3412 VSS.n5534 VSS.n5533 175.546
R3413 VSS.n5533 VSS.n35 175.546
R3414 VSS.n5529 VSS.n35 175.546
R3415 VSS.n5529 VSS.n37 175.546
R3416 VSS.n5525 VSS.n37 175.546
R3417 VSS.n5525 VSS.n40 175.546
R3418 VSS.n5521 VSS.n40 175.546
R3419 VSS.n5521 VSS.n42 175.546
R3420 VSS.n5517 VSS.n42 175.546
R3421 VSS.n5517 VSS.n44 175.546
R3422 VSS.n1136 VSS.n1133 175.546
R3423 VSS.n1140 VSS.n1133 175.546
R3424 VSS.n1140 VSS.n1130 175.546
R3425 VSS.n1159 VSS.n1130 175.546
R3426 VSS.n1159 VSS.n1131 175.546
R3427 VSS.n1155 VSS.n1131 175.546
R3428 VSS.n1155 VSS.n1144 175.546
R3429 VSS.n1151 VSS.n1144 175.546
R3430 VSS.n1151 VSS.n1148 175.546
R3431 VSS.n1148 VSS.n1146 175.546
R3432 VSS.n5500 VSS.n60 175.546
R3433 VSS.n5496 VSS.n60 175.546
R3434 VSS.n5496 VSS.n63 175.546
R3435 VSS.n5492 VSS.n63 175.546
R3436 VSS.n5492 VSS.n65 175.546
R3437 VSS.n5488 VSS.n65 175.546
R3438 VSS.n5488 VSS.n67 175.546
R3439 VSS.n5484 VSS.n67 175.546
R3440 VSS.n5484 VSS.n70 175.546
R3441 VSS.n5480 VSS.n70 175.546
R3442 VSS.n5480 VSS.n72 175.546
R3443 VSS.n4396 VSS.n4333 175.546
R3444 VSS.n4392 VSS.n4333 175.546
R3445 VSS.n4392 VSS.n4335 175.546
R3446 VSS.n4363 VSS.n4335 175.546
R3447 VSS.n4363 VSS.n4360 175.546
R3448 VSS.n4360 VSS.n4341 175.546
R3449 VSS.n4352 VSS.n4341 175.546
R3450 VSS.n4352 VSS.n4349 175.546
R3451 VSS.n4349 VSS.n336 175.546
R3452 VSS.n5292 VSS.n336 175.546
R3453 VSS.n5292 VSS.n337 175.546
R3454 VSS.n1523 VSS.n1491 175.546
R3455 VSS.n2559 VSS.n1491 175.546
R3456 VSS.n2559 VSS.n1492 175.546
R3457 VSS.n2555 VSS.n1492 175.546
R3458 VSS.n2555 VSS.n1527 175.546
R3459 VSS.n2548 VSS.n1527 175.546
R3460 VSS.n2548 VSS.n1534 175.546
R3461 VSS.n2544 VSS.n1534 175.546
R3462 VSS.n2544 VSS.n1536 175.546
R3463 VSS.n2537 VSS.n1536 175.546
R3464 VSS.n2537 VSS.n2535 175.546
R3465 VSS.n2528 VSS.n1563 175.546
R3466 VSS.n2524 VSS.n1563 175.546
R3467 VSS.n2524 VSS.n1565 175.546
R3468 VSS.n2235 VSS.n1565 175.546
R3469 VSS.n2235 VSS.n2230 175.546
R3470 VSS.n2244 VSS.n2230 175.546
R3471 VSS.n2247 VSS.n2244 175.546
R3472 VSS.n2247 VSS.n2225 175.546
R3473 VSS.n2285 VSS.n2225 175.546
R3474 VSS.n2285 VSS.n2223 175.546
R3475 VSS.n2289 VSS.n2223 175.546
R3476 VSS.n2298 VSS.n2296 175.546
R3477 VSS.n2298 VSS.n2127 175.546
R3478 VSS.n2309 VSS.n2127 175.546
R3479 VSS.n2309 VSS.n2125 175.546
R3480 VSS.n2313 VSS.n2125 175.546
R3481 VSS.n2315 VSS.n2313 175.546
R3482 VSS.n2315 VSS.n2120 175.546
R3483 VSS.n2326 VSS.n2120 175.546
R3484 VSS.n2326 VSS.n2118 175.546
R3485 VSS.n2330 VSS.n2118 175.546
R3486 VSS.n2330 VSS.n349 175.546
R3487 VSS.n5278 VSS.n5277 175.546
R3488 VSS.n5277 VSS.n351 175.546
R3489 VSS.n5273 VSS.n351 175.546
R3490 VSS.n5273 VSS.n354 175.546
R3491 VSS.n5269 VSS.n354 175.546
R3492 VSS.n5269 VSS.n357 175.546
R3493 VSS.n5265 VSS.n357 175.546
R3494 VSS.n5265 VSS.n359 175.546
R3495 VSS.n5261 VSS.n359 175.546
R3496 VSS.n5261 VSS.n361 175.546
R3497 VSS.n4966 VSS.n4963 175.546
R3498 VSS.n4966 VSS.n4961 175.546
R3499 VSS.n4971 VSS.n4961 175.546
R3500 VSS.n4971 VSS.n4958 175.546
R3501 VSS.n4975 VSS.n4958 175.546
R3502 VSS.n4976 VSS.n4975 175.546
R3503 VSS.n4979 VSS.n4976 175.546
R3504 VSS.n4979 VSS.n4956 175.546
R3505 VSS.n4984 VSS.n4956 175.546
R3506 VSS.n4984 VSS.n4953 175.546
R3507 VSS.n4989 VSS.n4953 175.546
R3508 VSS.n4992 VSS.n625 175.546
R3509 VSS.n4996 VSS.n625 175.546
R3510 VSS.n4996 VSS.n623 175.546
R3511 VSS.n5000 VSS.n623 175.546
R3512 VSS.n5000 VSS.n619 175.546
R3513 VSS.n5004 VSS.n619 175.546
R3514 VSS.n5004 VSS.n617 175.546
R3515 VSS.n5008 VSS.n617 175.546
R3516 VSS.n5008 VSS.n612 175.546
R3517 VSS.n5013 VSS.n612 175.546
R3518 VSS.n4654 VSS.n563 175.546
R3519 VSS.n5098 VSS.n563 175.546
R3520 VSS.n5098 VSS.n564 175.546
R3521 VSS.n5094 VSS.n564 175.546
R3522 VSS.n5094 VSS.n567 175.546
R3523 VSS.n572 VSS.n567 175.546
R3524 VSS.n5083 VSS.n572 175.546
R3525 VSS.n5083 VSS.n573 175.546
R3526 VSS.n5079 VSS.n573 175.546
R3527 VSS.n5079 VSS.n576 175.546
R3528 VSS.n5071 VSS.n576 175.546
R3529 VSS.n5043 VSS.n593 175.546
R3530 VSS.n5047 VSS.n593 175.546
R3531 VSS.n5047 VSS.n591 175.546
R3532 VSS.n5052 VSS.n591 175.546
R3533 VSS.n5052 VSS.n589 175.546
R3534 VSS.n5056 VSS.n589 175.546
R3535 VSS.n5056 VSS.n588 175.546
R3536 VSS.n5061 VSS.n588 175.546
R3537 VSS.n5061 VSS.n586 175.546
R3538 VSS.n5065 VSS.n586 175.546
R3539 VSS.n5067 VSS.n5065 175.546
R3540 VSS.n5018 VSS.n606 175.546
R3541 VSS.n5018 VSS.n604 175.546
R3542 VSS.n5023 VSS.n604 175.546
R3543 VSS.n5023 VSS.n602 175.546
R3544 VSS.n5027 VSS.n602 175.546
R3545 VSS.n5027 VSS.n601 175.546
R3546 VSS.n5031 VSS.n601 175.546
R3547 VSS.n5031 VSS.n599 175.546
R3548 VSS.n5036 VSS.n599 175.546
R3549 VSS.n5036 VSS.n595 175.546
R3550 VSS.n5254 VSS.n366 175.546
R3551 VSS.n5250 VSS.n366 175.546
R3552 VSS.n5250 VSS.n369 175.546
R3553 VSS.n5246 VSS.n369 175.546
R3554 VSS.n5246 VSS.n372 175.546
R3555 VSS.n5242 VSS.n372 175.546
R3556 VSS.n5242 VSS.n376 175.546
R3557 VSS.n5238 VSS.n376 175.546
R3558 VSS.n5238 VSS.n378 175.546
R3559 VSS.n5234 VSS.n378 175.546
R3560 VSS.n4426 VSS.n894 175.546
R3561 VSS.n4529 VSS.n894 175.546
R3562 VSS.n4529 VSS.n895 175.546
R3563 VSS.n4525 VSS.n895 175.546
R3564 VSS.n4525 VSS.n4430 175.546
R3565 VSS.n4435 VSS.n4430 175.546
R3566 VSS.n4514 VSS.n4435 175.546
R3567 VSS.n4514 VSS.n4436 175.546
R3568 VSS.n4510 VSS.n4436 175.546
R3569 VSS.n4510 VSS.n4439 175.546
R3570 VSS.n4502 VSS.n4439 175.546
R3571 VSS.n4605 VSS.n781 175.546
R3572 VSS.n4635 VSS.n781 175.546
R3573 VSS.n4635 VSS.n782 175.546
R3574 VSS.n4631 VSS.n782 175.546
R3575 VSS.n4631 VSS.n4609 175.546
R3576 VSS.n4617 VSS.n4609 175.546
R3577 VSS.n4620 VSS.n4617 175.546
R3578 VSS.n4620 VSS.n739 175.546
R3579 VSS.n4645 VSS.n739 175.546
R3580 VSS.n4645 VSS.n735 175.546
R3581 VSS.n4650 VSS.n735 175.546
R3582 VSS.n3724 VSS.n3721 175.546
R3583 VSS.n3728 VSS.n3721 175.546
R3584 VSS.n3728 VSS.n3719 175.546
R3585 VSS.n3732 VSS.n3719 175.546
R3586 VSS.n3732 VSS.n3717 175.546
R3587 VSS.n3737 VSS.n3717 175.546
R3588 VSS.n3737 VSS.n3715 175.546
R3589 VSS.n3742 VSS.n3715 175.546
R3590 VSS.n3742 VSS.n3714 175.546
R3591 VSS.n3746 VSS.n3714 175.546
R3592 VSS.n3747 VSS.n3746 175.546
R3593 VSS.n3754 VSS.n1194 175.546
R3594 VSS.n4004 VSS.n1194 175.546
R3595 VSS.n4004 VSS.n1195 175.546
R3596 VSS.n4000 VSS.n1195 175.546
R3597 VSS.n4000 VSS.n1198 175.546
R3598 VSS.n1205 VSS.n1198 175.546
R3599 VSS.n1209 VSS.n1204 175.546
R3600 VSS.n1214 VSS.n1213 175.546
R3601 VSS.n3989 VSS.n1201 175.546
R3602 VSS.n3989 VSS.n1218 175.546
R3603 VSS.n3985 VSS.n1218 175.546
R3604 VSS.n3985 VSS.n1221 175.546
R3605 VSS.n1230 VSS.n1221 175.546
R3606 VSS.n3976 VSS.n1230 175.546
R3607 VSS.n3976 VSS.n1231 175.546
R3608 VSS.n3972 VSS.n1231 175.546
R3609 VSS.n3972 VSS.n1233 175.546
R3610 VSS.n3964 VSS.n1233 175.546
R3611 VSS.n3964 VSS.n1242 175.546
R3612 VSS.n3957 VSS.n1273 175.546
R3613 VSS.n3941 VSS.n1273 175.546
R3614 VSS.n3941 VSS.n1281 175.546
R3615 VSS.n3946 VSS.n1281 175.546
R3616 VSS.n3946 VSS.n3940 175.546
R3617 VSS.n3940 VSS.n1282 175.546
R3618 VSS.n1289 VSS.n1282 175.546
R3619 VSS.n3931 VSS.n1289 175.546
R3620 VSS.n3931 VSS.n1290 175.546
R3621 VSS.n3927 VSS.n1290 175.546
R3622 VSS.n3927 VSS.n1294 175.546
R3623 VSS.t18 VSS.n340 173.071
R3624 VSS.n5258 VSS.t72 170.631
R3625 VSS.n4987 VSS.t72 170.631
R3626 VSS.n5011 VSS.t72 170.631
R3627 VSS.n5039 VSS.t72 170.631
R3628 VSS.n341 VSS.t104 164.196
R3629 VSS.n1167 VSS.n1166 159.255
R3630 VSS.n3994 VSS.n1202 152.643
R3631 VSS.n4281 VSS.n1042 150
R3632 VSS.n4289 VSS.n4288 150
R3633 VSS.n4297 VSS.n4296 150
R3634 VSS.n4312 VSS.n4165 150
R3635 VSS.n4124 VSS.n4123 150
R3636 VSS.n4128 VSS.n4127 150
R3637 VSS.n4132 VSS.n4131 150
R3638 VSS.n4136 VSS.n4135 150
R3639 VSS.n4139 VSS.n1055 150
R3640 VSS.n4158 VSS.n1056 150
R3641 VSS.n1086 VSS.n1085 150
R3642 VSS.n1076 VSS.n1075 150
R3643 VSS.n4164 VSS.n4160 150
R3644 VSS.n4177 VSS.n4160 150
R3645 VSS.n4175 VSS.n4174 150
R3646 VSS.n4171 VSS.n4170 150
R3647 VSS.n4167 VSS.n1051 150
R3648 VSS.n5468 VSS.n86 150
R3649 VSS.n5466 VSS.n87 150
R3650 VSS.n133 VSS.n132 150
R3651 VSS.n5449 VSS.n140 150
R3652 VSS.n5432 VSS.n145 150
R3653 VSS.n5436 VSS.n5434 150
R3654 VSS.n5440 VSS.n143 150
R3655 VSS.n5443 VSS.n5442 150
R3656 VSS.n4153 VSS.n1060 150
R3657 VSS.n4155 VSS.n1059 150
R3658 VSS.n1094 VSS.n1071 150
R3659 VSS.n1097 VSS.n1096 150
R3660 VSS.n4062 VSS.n4060 150
R3661 VSS.n4058 VSS.n1109 150
R3662 VSS.n4054 VSS.n4052 150
R3663 VSS.n4052 VSS.n4051 150
R3664 VSS.n4049 VSS.n1113 150
R3665 VSS.n5463 VSS.n91 150
R3666 VSS.n129 VSS.n92 150
R3667 VSS.n137 VSS.n136 150
R3668 VSS.n5460 VSS.n111 150
R3669 VSS.n4039 VSS.n4038 150
R3670 VSS.n4035 VSS.n4034 150
R3671 VSS.n4031 VSS.n4030 150
R3672 VSS.n4027 VSS.n4026 150
R3673 VSS.n3780 VSS.n3779 150
R3674 VSS.n3791 VSS.n3790 150
R3675 VSS.n3557 VSS.n3556 150
R3676 VSS.n3570 VSS.n3569 150
R3677 VSS.n110 VSS.n106 150
R3678 VSS.n3509 VSS.n106 150
R3679 VSS.n3513 VSS.n3512 150
R3680 VSS.n3517 VSS.n3516 150
R3681 VSS.n3519 VSS.n101 150
R3682 VSS.n3651 VSS.n3650 150
R3683 VSS.n3660 VSS.n3659 150
R3684 VSS.n3669 VSS.n3668 150
R3685 VSS.n3679 VSS.n3678 150
R3686 VSS.n3591 VSS.n3548 150
R3687 VSS.n3595 VSS.n3594 150
R3688 VSS.n3599 VSS.n3598 150
R3689 VSS.n3603 VSS.n3602 150
R3690 VSS.n3784 VSS.n3778 150
R3691 VSS.n3787 VSS.n3533 150
R3692 VSS.n3575 VSS.n3534 150
R3693 VSS.n3566 VSS.n3551 150
R3694 VSS.n3777 VSS.n3776 150
R3695 VSS.n3773 VSS.n3772 150
R3696 VSS.n3769 VSS.n3543 150
R3697 VSS.n3766 VSS.n3543 150
R3698 VSS.n3764 VSS.n3763 150
R3699 VSS.n3648 VSS.n3647 150
R3700 VSS.n3645 VSS.n3644 150
R3701 VSS.n3642 VSS.n3641 150
R3702 VSS.n3682 VSS.n3610 150
R3703 VSS.n3638 VSS.n3637 150
R3704 VSS.n3637 VSS.n3617 150
R3705 VSS.n3633 VSS.n3632 150
R3706 VSS.n3630 VSS.n3620 150
R3707 VSS.n3626 VSS.n3625 150
R3708 VSS.n3623 VSS.n3622 150
R3709 VSS.n3982 VSS.n3981 150
R3710 VSS.n3979 VSS.n1227 150
R3711 VSS.n3969 VSS.n1239 150
R3712 VSS.n3703 VSS.n3702 150
R3713 VSS.n3700 VSS.n3685 150
R3714 VSS.n3696 VSS.n3695 150
R3715 VSS.n3693 VSS.n3689 150
R3716 VSS.n3476 VSS.n3475 150
R3717 VSS.n3462 VSS.n3460 150
R3718 VSS.n3464 VSS.n3459 150
R3719 VSS.n3873 VSS.n1307 150
R3720 VSS.n3444 VSS.n3424 150
R3721 VSS.n3440 VSS.n3424 150
R3722 VSS.n3438 VSS.n3437 150
R3723 VSS.n3435 VSS.n3428 150
R3724 VSS.n3431 VSS.n3430 150
R3725 VSS.n3952 VSS.n3951 150
R3726 VSS.n3949 VSS.n1278 150
R3727 VSS.n3937 VSS.n3936 150
R3728 VSS.n3934 VSS.n1286 150
R3729 VSS.n3878 VSS.n3876 150
R3730 VSS.n3882 VSS.n1302 150
R3731 VSS.n3885 VSS.n3884 150
R3732 VSS.n3889 VSS.n3888 150
R3733 VSS.n5101 VSS.n560 150
R3734 VSS.n5091 VSS.n5090 150
R3735 VSS.n5087 VSS.n5086 150
R3736 VSS.n579 VSS.n578 150
R3737 VSS.n4706 VSS.n4705 150
R3738 VSS.n4702 VSS.n4701 150
R3739 VSS.n4698 VSS.n4697 150
R3740 VSS.n4694 VSS.n4693 150
R3741 VSS.n4744 VSS.n541 150
R3742 VSS.n4752 VSS.n4751 150
R3743 VSS.n4760 VSS.n4759 150
R3744 VSS.n4767 VSS.n4766 150
R3745 VSS.n721 VSS.n548 150
R3746 VSS.n724 VSS.n548 150
R3747 VSS.n728 VSS.n727 150
R3748 VSS.n730 VSS.n553 150
R3749 VSS.n559 VSS.n553 150
R3750 VSS.n5107 VSS.n537 150
R3751 VSS.n4748 VSS.n4747 150
R3752 VSS.n4756 VSS.n4755 150
R3753 VSS.n4764 VSS.n4763 150
R3754 VSS.n4710 VSS.n4709 150
R3755 VSS.n4714 VSS.n4713 150
R3756 VSS.n4718 VSS.n4717 150
R3757 VSS.n4722 VSS.n4721 150
R3758 VSS.n5110 VSS.n517 150
R3759 VSS.n4842 VSS.n518 150
R3760 VSS.n4866 VSS.n4865 150
R3761 VSS.n4875 VSS.n4874 150
R3762 VSS.n4795 VSS.n525 150
R3763 VSS.n4792 VSS.n525 150
R3764 VSS.n4790 VSS.n4789 150
R3765 VSS.n4786 VSS.n530 150
R3766 VSS.n536 VSS.n530 150
R3767 VSS.n4935 VSS.n4934 150
R3768 VSS.n4923 VSS.n4827 150
R3769 VSS.n4921 VSS.n4828 150
R3770 VSS.n4902 VSS.n4900 150
R3771 VSS.n4820 VSS.n663 150
R3772 VSS.n4816 VSS.n663 150
R3773 VSS.n4814 VSS.n4813 150
R3774 VSS.n4811 VSS.n667 150
R3775 VSS.n4807 VSS.n4806 150
R3776 VSS.n5115 VSS.n512 150
R3777 VSS.n5113 VSS.n513 150
R3778 VSS.n4857 VSS.n4852 150
R3779 VSS.n4855 VSS.n4854 150
R3780 VSS.n4897 VSS.n4830 150
R3781 VSS.n4893 VSS.n4892 150
R3782 VSS.n4890 VSS.n4835 150
R3783 VSS.n4886 VSS.n4885 150
R3784 VSS.n5158 VSS.n446 150
R3785 VSS.n463 VSS.n461 150
R3786 VSS.n5144 VSS.n5143 150
R3787 VSS.n5141 VSS.n466 150
R3788 VSS.n1865 VSS.n1864 150
R3789 VSS.n1862 VSS.n1844 150
R3790 VSS.n1858 VSS.n1857 150
R3791 VSS.n1855 VSS.n1847 150
R3792 VSS.n5177 VSS.n5176 150
R3793 VSS.n5179 VSS.n436 150
R3794 VSS.n1840 VSS.n1819 150
R3795 VSS.n1868 VSS.n1842 150
R3796 VSS.n5174 VSS.n437 150
R3797 VSS.n5170 VSS.n5169 150
R3798 VSS.n5167 VSS.n443 150
R3799 VSS.n5163 VSS.n443 150
R3800 VSS.n5161 VSS.n5160 150
R3801 VSS.n789 VSS.n788 150
R3802 VSS.n4579 VSS.n4578 150
R3803 VSS.n807 VSS.n806 150
R3804 VSS.n4566 VSS.n4565 150
R3805 VSS.n816 VSS.n483 150
R3806 VSS.n820 VSS.n819 150
R3807 VSS.n824 VSS.n823 150
R3808 VSS.n828 VSS.n827 150
R3809 VSS.n5155 VSS.n5154 150
R3810 VSS.n5132 VSS.n5131 150
R3811 VSS.n5136 VSS.n5134 150
R3812 VSS.n5138 VSS.n469 150
R3813 VSS.n3175 VSS.n3174 150
R3814 VSS.n3171 VSS.n3170 150
R3815 VSS.n3167 VSS.n478 150
R3816 VSS.n3164 VSS.n478 150
R3817 VSS.n3162 VSS.n3161 150
R3818 VSS.n4638 VSS.n778 150
R3819 VSS.n4628 VSS.n4627 150
R3820 VSS.n4624 VSS.n4623 150
R3821 VSS.n4615 VSS.n4614 150
R3822 VSS.n760 VSS.n759 150
R3823 VSS.n764 VSS.n763 150
R3824 VSS.n766 VSS.n757 150
R3825 VSS.n771 VSS.n745 150
R3826 VSS.n796 VSS.n795 150
R3827 VSS.n4575 VSS.n4574 150
R3828 VSS.n811 VSS.n810 150
R3829 VSS.n4562 VSS.n4561 150
R3830 VSS.n4590 VSS.n753 150
R3831 VSS.n4593 VSS.n753 150
R3832 VSS.n4597 VSS.n4596 150
R3833 VSS.n4599 VSS.n773 150
R3834 VSS.n777 VSS.n773 150
R3835 VSS.n4532 VSS.n891 150
R3836 VSS.n4522 VSS.n4521 150
R3837 VSS.n4518 VSS.n4517 150
R3838 VSS.n4442 VSS.n4441 150
R3839 VSS.n4449 VSS.n4448 150
R3840 VSS.n4453 VSS.n4452 150
R3841 VSS.n4457 VSS.n4456 150
R3842 VSS.n4461 VSS.n4460 150
R3843 VSS.n907 VSS.n870 150
R3844 VSS.n935 VSS.n934 150
R3845 VSS.n920 VSS.n919 150
R3846 VSS.n873 VSS.n872 150
R3847 VSS.n4411 VSS.n879 150
R3848 VSS.n4414 VSS.n879 150
R3849 VSS.n4418 VSS.n4417 150
R3850 VSS.n4420 VSS.n884 150
R3851 VSS.n890 VSS.n884 150
R3852 VSS.n2428 VSS.n2427 150
R3853 VSS.n2425 VSS.n2037 150
R3854 VSS.n2413 VSS.n2412 150
R3855 VSS.n2410 VSS.n2050 150
R3856 VSS.n2364 VSS.n2066 150
R3857 VSS.n2368 VSS.n2366 150
R3858 VSS.n2372 VSS.n2064 150
R3859 VSS.n2375 VSS.n2374 150
R3860 VSS.n2450 VSS.n2449 150
R3861 VSS.n2452 VSS.n2012 150
R3862 VSS.n2102 VSS.n2083 150
R3863 VSS.n2104 VSS.n2081 150
R3864 VSS.n2447 VSS.n2446 150
R3865 VSS.n2444 VSS.n2014 150
R3866 VSS.n2440 VSS.n2438 150
R3867 VSS.n2438 VSS.n2437 150
R3868 VSS.n2435 VSS.n2017 150
R3869 VSS.n4938 VSS.n657 150
R3870 VSS.n4926 VSS.n4925 150
R3871 VSS.n4914 VSS.n4913 150
R3872 VSS.n4907 VSS.n4906 150
R3873 VSS.n2390 VSS.n2389 150
R3874 VSS.n2386 VSS.n2385 150
R3875 VSS.n2382 VSS.n2381 150
R3876 VSS.n2378 VSS.n639 150
R3877 VSS.n2422 VSS.n2421 150
R3878 VSS.n2046 VSS.n2045 150
R3879 VSS.n2407 VSS.n2406 150
R3880 VSS.n2059 VSS.n2058 150
R3881 VSS.n2029 VSS.n647 150
R3882 VSS.n2026 VSS.n647 150
R3883 VSS.n2024 VSS.n2023 150
R3884 VSS.n2020 VSS.n652 150
R3885 VSS.n656 VSS.n652 150
R3886 VSS.n2457 VSS.n2008 150
R3887 VSS.n2455 VSS.n2009 150
R3888 VSS.n2096 VSS.n2094 150
R3889 VSS.n2108 VSS.n2077 150
R3890 VSS.n2337 VSS.n2335 150
R3891 VSS.n2341 VSS.n2112 150
R3892 VSS.n2345 VSS.n2343 150
R3893 VSS.n2349 VSS.n2110 150
R3894 VSS.n2306 VSS.n2304 150
R3895 VSS.n2318 VSS.n2123 150
R3896 VSS.n2322 VSS.n2320 150
R3897 VSS.n2333 VSS.n2114 150
R3898 VSS.n2149 VSS.n2147 150
R3899 VSS.n2147 VSS.n2146 150
R3900 VSS.n2143 VSS.n2142 150
R3901 VSS.n2140 VSS.n2137 150
R3902 VSS.n2137 VSS.n2136 150
R3903 VSS.n2501 VSS.n1576 150
R3904 VSS.n2489 VSS.n1589 150
R3905 VSS.n2487 VSS.n1590 150
R3906 VSS.n2260 VSS.n2259 150
R3907 VSS.n2280 VSS.n2254 150
R3908 VSS.n2276 VSS.n2274 150
R3909 VSS.n2272 VSS.n2256 150
R3910 VSS.n2268 VSS.n2266 150
R3911 VSS.n2521 VSS.n1569 150
R3912 VSS.n2241 VSS.n2239 150
R3913 VSS.n2251 VSS.n2228 150
R3914 VSS.n2282 VSS.n2253 150
R3915 VSS.n2515 VSS.n2514 150
R3916 VSS.n2514 VSS.n2513 150
R3917 VSS.n2510 VSS.n2509 150
R3918 VSS.n2507 VSS.n1574 150
R3919 VSS.n2503 VSS.n1574 150
R3920 VSS.n3043 VSS.n1484 150
R3921 VSS.n3006 VSS.n3005 150
R3922 VSS.n3029 VSS.n3028 150
R3923 VSS.n3019 VSS.n3018 150
R3924 VSS.n1555 VSS.n1554 150
R3925 VSS.n1551 VSS.n1550 150
R3926 VSS.n1547 VSS.n1546 150
R3927 VSS.n1543 VSS.n1466 150
R3928 VSS.n1530 VSS.n1529 150
R3929 VSS.n2552 VSS.n2551 150
R3930 VSS.n1539 VSS.n1538 150
R3931 VSS.n2541 VSS.n2540 150
R3932 VSS.n2565 VSS.n1474 150
R3933 VSS.n2568 VSS.n1474 150
R3934 VSS.n2572 VSS.n2571 150
R3935 VSS.n2574 VSS.n1479 150
R3936 VSS.n1483 VSS.n1479 150
R3937 VSS.n5357 VSS.n5356 150
R3938 VSS.n5354 VSS.n310 150
R3939 VSS.n2685 VSS.n2680 150
R3940 VSS.n2690 VSS.n2689 150
R3941 VSS.n5299 VSS.n5297 150
R3942 VSS.n5303 VSS.n331 150
R3943 VSS.n5307 VSS.n5305 150
R3944 VSS.n5311 VSS.n329 150
R3945 VSS.n4389 VSS.n4366 150
R3946 VSS.n4357 VSS.n4343 150
R3947 VSS.n4355 VSS.n4345 150
R3948 VSS.n5295 VSS.n333 150
R3949 VSS.n4383 VSS.n4382 150
R3950 VSS.n4382 VSS.n4381 150
R3951 VSS.n4378 VSS.n4377 150
R3952 VSS.n4375 VSS.n4372 150
R3953 VSS.n4372 VSS.n4371 150
R3954 VSS.n4076 VSS.n4075 150
R3955 VSS.n4093 VSS.n4092 150
R3956 VSS.n4082 VSS.n4081 150
R3957 VSS.n4321 VSS.n1018 150
R3958 VSS.n4106 VSS.n1026 150
R3959 VSS.n4109 VSS.n1026 150
R3960 VSS.n4113 VSS.n4112 150
R3961 VSS.n4115 VSS.n1031 150
R3962 VSS.n1037 VSS.n1031 150
R3963 VSS.n4318 VSS.n1038 150
R3964 VSS.n4285 VSS.n4284 150
R3965 VSS.n4293 VSS.n4292 150
R3966 VSS.n4301 VSS.n4300 150
R3967 VSS.n4182 VSS.n1019 150
R3968 VSS.n4186 VSS.n4185 150
R3969 VSS.n4190 VSS.n4189 150
R3970 VSS.n4194 VSS.n4193 150
R3971 VSS.n1769 VSS.n1768 150
R3972 VSS.n1776 VSS.n1775 150
R3973 VSS.n1789 VSS.n1788 150
R3974 VSS.n1710 VSS.n1709 150
R3975 VSS.n1994 VSS.n1607 150
R3976 VSS.n1992 VSS.n1991 150
R3977 VSS.n1988 VSS.n1987 150
R3978 VSS.n1984 VSS.n1983 150
R3979 VSS.n2498 VSS.n2497 150
R3980 VSS.n2482 VSS.n2481 150
R3981 VSS.n2484 VSS.n1593 150
R3982 VSS.n2479 VSS.n1609 150
R3983 VSS.n1727 VSS.n1726 150
R3984 VSS.n1731 VSS.n1730 150
R3985 VSS.n1733 VSS.n1602 150
R3986 VSS.n1736 VSS.n1602 150
R3987 VSS.n1740 VSS.n1739 150
R3988 VSS.n5184 VSS.n431 150
R3989 VSS.n5182 VSS.n432 150
R3990 VSS.n1831 VSS.n1821 150
R3991 VSS.n1835 VSS.n1834 150
R3992 VSS.n1974 VSS.n1804 150
R3993 VSS.n1970 VSS.n1968 150
R3994 VSS.n1966 VSS.n1806 150
R3995 VSS.n1962 VSS.n1960 150
R3996 VSS.n1781 VSS.n1719 150
R3997 VSS.n1785 VSS.n1783 150
R3998 VSS.n1801 VSS.n1707 150
R3999 VSS.n1976 VSS.n1803 150
R4000 VSS.n1760 VSS.n1759 150
R4001 VSS.n1759 VSS.n1758 150
R4002 VSS.n1755 VSS.n1754 150
R4003 VSS.n1752 VSS.n1746 150
R4004 VSS.n1748 VSS.n1746 150
R4005 VSS.n2970 VSS.n2584 150
R4006 VSS.n2939 VSS.n2935 150
R4007 VSS.n2955 VSS.n2954 150
R4008 VSS.n3076 VSS.n1450 150
R4009 VSS.n3059 VSS.n1455 150
R4010 VSS.n3063 VSS.n3061 150
R4011 VSS.n3067 VSS.n1453 150
R4012 VSS.n3070 VSS.n3069 150
R4013 VSS.n3040 VSS.n3039 150
R4014 VSS.n3011 VSS.n3010 150
R4015 VSS.n3025 VSS.n3013 150
R4016 VSS.n3023 VSS.n3016 150
R4017 VSS.n2986 VSS.n1487 150
R4018 VSS.n2982 VSS.n2981 150
R4019 VSS.n2979 VSS.n2581 150
R4020 VSS.n2975 VSS.n2581 150
R4021 VSS.n2973 VSS.n2972 150
R4022 VSS.n2850 VSS.n2734 150
R4023 VSS.n2831 VSS.n2821 150
R4024 VSS.n2836 VSS.n2835 150
R4025 VSS.n3109 VSS.n3108 150
R4026 VSS.n3091 VSS.n3089 150
R4027 VSS.n3095 VSS.n1439 150
R4028 VSS.n3099 VSS.n3097 150
R4029 VSS.n3103 VSS.n1437 150
R4030 VSS.n2965 VSS.n2588 150
R4031 VSS.n2948 VSS.n2947 150
R4032 VSS.n2950 VSS.n2945 150
R4033 VSS.n3087 VSS.n1441 150
R4034 VSS.n2865 VSS.n2863 150
R4035 VSS.n2863 VSS.n2862 150
R4036 VSS.n2859 VSS.n2858 150
R4037 VSS.n2856 VSS.n2731 150
R4038 VSS.n2852 VSS.n2731 150
R4039 VSS.n5420 VSS.n165 150
R4040 VSS.n5418 VSS.n166 150
R4041 VSS.n2661 VSS.n2659 150
R4042 VSS.n2671 VSS.n2647 150
R4043 VSS.n2703 VSS.n2701 150
R4044 VSS.n2707 VSS.n2675 150
R4045 VSS.n2711 VSS.n2709 150
R4046 VSS.n2715 VSS.n2673 150
R4047 VSS.n5349 VSS.n5347 150
R4048 VSS.n5351 VSS.n5324 150
R4049 VSS.n2695 VSS.n2678 150
R4050 VSS.n2698 VSS.n2697 150
R4051 VSS.n5345 VSS.n5344 150
R4052 VSS.n5342 VSS.n5326 150
R4053 VSS.n5338 VSS.n5336 150
R4054 VSS.n5336 VSS.n5335 150
R4055 VSS.n5333 VSS.n5330 150
R4056 VSS.n5412 VSS.n190 150
R4057 VSS.n5400 VSS.n5399 150
R4058 VSS.n226 VSS.n225 150
R4059 VSS.n5386 VSS.n5385 150
R4060 VSS.n2637 VSS.n2636 150
R4061 VSS.n2633 VSS.n2632 150
R4062 VSS.n2629 VSS.n2628 150
R4063 VSS.n2625 VSS.n2624 150
R4064 VSS.n5415 VSS.n170 150
R4065 VSS.n2656 VSS.n171 150
R4066 VSS.n2667 VSS.n2666 150
R4067 VSS.n2645 VSS.n2644 150
R4068 VSS.n3268 VSS.n178 150
R4069 VSS.n3271 VSS.n178 150
R4070 VSS.n3275 VSS.n3274 150
R4071 VSS.n3277 VSS.n183 150
R4072 VSS.n189 VSS.n183 150
R4073 VSS.n2792 VSS.n2743 150
R4074 VSS.n2763 VSS.n2751 150
R4075 VSS.n2761 VSS.n2752 150
R4076 VSS.n3144 VSS.n3143 150
R4077 VSS.n3126 VSS.n3124 150
R4078 VSS.n3130 VSS.n1419 150
R4079 VSS.n3134 VSS.n3132 150
R4080 VSS.n3138 VSS.n1417 150
R4081 VSS.n2847 VSS.n2846 150
R4082 VSS.n2827 VSS.n2826 150
R4083 VSS.n2824 VSS.n2823 150
R4084 VSS.n3121 VSS.n1422 150
R4085 VSS.n2808 VSS.n2737 150
R4086 VSS.n2804 VSS.n2803 150
R4087 VSS.n2801 VSS.n2740 150
R4088 VSS.n2797 VSS.n2740 150
R4089 VSS.n2795 VSS.n2794 150
R4090 VSS.n4538 VSS.n866 150
R4091 VSS.n939 VSS.n938 150
R4092 VSS.n916 VSS.n915 150
R4093 VSS.n925 VSS.n924 150
R4094 VSS.n1403 VSS.n1402 150
R4095 VSS.n1399 VSS.n1398 150
R4096 VSS.n1395 VSS.n1394 150
R4097 VSS.n1391 VSS.n848 150
R4098 VSS.n2769 VSS.n2768 150
R4099 VSS.n2758 VSS.n2757 150
R4100 VSS.n1414 VSS.n1413 150
R4101 VSS.n3155 VSS.n3154 150
R4102 VSS.n2785 VSS.n856 150
R4103 VSS.n2782 VSS.n856 150
R4104 VSS.n2780 VSS.n2779 150
R4105 VSS.n2776 VSS.n861 150
R4106 VSS.n865 VSS.n861 150
R4107 VSS.n3502 VSS.n3501 150
R4108 VSS.n3376 VSS.n3375 150
R4109 VSS.n3405 VSS.n3404 150
R4110 VSS.n3388 VSS.n3387 150
R4111 VSS.n1325 VSS.n217 150
R4112 VSS.n1329 VSS.n1328 150
R4113 VSS.n1333 VSS.n1332 150
R4114 VSS.n1337 VSS.n1336 150
R4115 VSS.n5409 VSS.n5408 150
R4116 VSS.n5397 VSS.n202 150
R4117 VSS.n5394 VSS.n203 150
R4118 VSS.n5383 VSS.n219 150
R4119 VSS.n3352 VSS.n3351 150
R4120 VSS.n3356 VSS.n3355 150
R4121 VSS.n3358 VSS.n212 150
R4122 VSS.n3361 VSS.n212 150
R4123 VSS.n3365 VSS.n3364 150
R4124 VSS.n3479 VSS.n3419 150
R4125 VSS.n3470 VSS.n3469 150
R4126 VSS.n3467 VSS.n3453 150
R4127 VSS.n3863 VSS.n3862 150
R4128 VSS.n3845 VSS.n3843 150
R4129 VSS.n3849 VSS.n1321 150
R4130 VSS.n3853 VSS.n3851 150
R4131 VSS.n3857 VSS.n1319 150
R4132 VSS.n3498 VSS.n3413 150
R4133 VSS.n3399 VSS.n3398 150
R4134 VSS.n3401 VSS.n3397 150
R4135 VSS.n3841 VSS.n1323 150
R4136 VSS.n3493 VSS.n3414 150
R4137 VSS.n3489 VSS.n3414 150
R4138 VSS.n3487 VSS.n3486 150
R4139 VSS.n3483 VSS.n3482 150
R4140 VSS.n3482 VSS.n3481 150
R4141 VSS.n1191 VSS.n1190 146.299
R4142 VSS.n3995 VSS.n1201 146.287
R4143 VSS.t72 VSS.n353 138.78
R4144 VSS.n5245 VSS.t72 138.78
R4145 VSS.n4974 VSS.t72 138.78
R4146 VSS.t72 VSS.n5001 138.78
R4147 VSS.n5021 VSS.t72 138.78
R4148 VSS.n5050 VSS.t72 138.78
R4149 VSS.n5071 VSS.n584 138.486
R4150 VSS.n1695 VSS.t57 130.675
R4151 VSS.n1795 VSS.t57 130.675
R4152 VSS.n1874 VSS.t57 130.675
R4153 VSS.n454 VSS.t57 130.675
R4154 VSS.n4555 VSS.t57 130.675
R4155 VSS.n3149 VSS.t69 130.675
R4156 VSS.n5319 VSS.t60 130.675
R4157 VSS.n2723 VSS.t60 130.675
R4158 VSS.n3342 VSS.t60 130.675
R4159 VSS.n1344 VSS.t60 130.675
R4160 VSS.n3868 VSS.t60 130.675
R4161 VSS.n2467 VSS.n1999 129.708
R4162 VSS.n1926 VSS.n389 129.708
R4163 VSS.n1919 VSS.n1918 129.708
R4164 VSS.n681 VSS.n499 129.708
R4165 VSS.n4683 VSS.n4682 129.708
R4166 VSS.n5371 VSS.n291 129.708
R4167 VSS.n2923 VSS.n2593 129.708
R4168 VSS.n5374 VSS.n5373 129.708
R4169 VSS.n3254 VSS.n1346 129.708
R4170 VSS.n950 VSS.n949 129.708
R4171 VSS.n1650 VSS.n1460 129.708
R4172 VSS.n5221 VSS.n400 129.708
R4173 VSS.n5193 VSS.n5191 129.708
R4174 VSS.n3215 VSS.n1388 129.708
R4175 VSS.n4470 VSS.n837 129.708
R4176 VSS.n970 VSS.n302 129.708
R4177 VSS.n1007 VSS.n152 129.708
R4178 VSS.n3341 VSS.n983 129.708
R4179 VSS.n3831 VSS.n3261 129.708
R4180 VSS.n4401 VSS.n956 129.708
R4181 VSS.n1584 VSS.t57 128.062
R4182 VSS.n5225 VSS.t57 128.062
R4183 VSS.n5189 VSS.t57 128.062
R4184 VSS.n456 VSS.t57 128.062
R4185 VSS.n792 VSS.t57 128.062
R4186 VSS.n3223 VSS.t69 128.062
R4187 VSS.n5364 VSS.t60 128.062
R4188 VSS.n5425 VSS.t60 128.062
R4189 VSS.n198 VSS.t60 128.062
R4190 VSS.n3835 VSS.t60 128.062
R4191 VSS.n4405 VSS.t60 128.062
R4192 VSS.n5538 VSS.n29 124.832
R4193 VSS.n46 VSS.n44 124.832
R4194 VSS.n1146 VSS.n1125 124.832
R4195 VSS.n5475 VSS.n72 124.832
R4196 VSS.n363 VSS.n361 124.832
R4197 VSS.n4989 VSS.n4954 124.832
R4198 VSS.n5013 VSS.n615 124.832
R4199 VSS.n5041 VSS.n595 124.832
R4200 VSS.n5234 VSS.n380 124.832
R4201 VSS.n3747 VSS.n3583 124.832
R4202 VSS.n1168 VSS.n339 119.819
R4203 VSS.n3996 VSS.n1200 113.022
R4204 VSS.n3959 VSS.n3958 113.022
R4205 VSS.n4427 VSS.n896 113.022
R4206 VSS.n4606 VSS.n783 113.022
R4207 VSS.n4653 VSS.n4652 113.022
R4208 VSS.n3962 VSS.n3961 107.427
R4209 VSS.n3893 VSS.n1293 107.427
R4210 VSS.n4501 VSS.n4500 107.427
R4211 VSS.n4649 VSS.n4648 107.427
R4212 VSS.n5070 VSS.n5069 107.427
R4213 VSS.n3988 VSS.n3987 100.713
R4214 VSS.n3987 VSS.n3986 100.713
R4215 VSS.n3986 VSS.n1220 100.713
R4216 VSS.n1229 VSS.n1220 100.713
R4217 VSS.n3975 VSS.n3974 100.713
R4218 VSS.n3974 VSS.n3973 100.713
R4219 VSS.n3973 VSS.n1232 100.713
R4220 VSS.n3963 VSS.n1232 100.713
R4221 VSS.n3963 VSS.n3962 100.713
R4222 VSS.n3958 VSS.n1272 100.713
R4223 VSS.n3942 VSS.n1272 100.713
R4224 VSS.n3943 VSS.n3942 100.713
R4225 VSS.n3945 VSS.n3943 100.713
R4226 VSS.n3945 VSS.n3944 100.713
R4227 VSS.n1292 VSS.n1291 100.713
R4228 VSS.n3930 VSS.n1292 100.713
R4229 VSS.n3930 VSS.n3929 100.713
R4230 VSS.n3929 VSS.n3928 100.713
R4231 VSS.n3928 VSS.n1293 100.713
R4232 VSS.n4428 VSS.n4427 100.713
R4233 VSS.n4528 VSS.n4428 100.713
R4234 VSS.n4528 VSS.n4527 100.713
R4235 VSS.n4527 VSS.n4526 100.713
R4236 VSS.n4526 VSS.n4429 100.713
R4237 VSS.n4513 VSS.n4437 100.713
R4238 VSS.n4513 VSS.n4512 100.713
R4239 VSS.n4512 VSS.n4511 100.713
R4240 VSS.n4511 VSS.n4438 100.713
R4241 VSS.n4501 VSS.n4438 100.713
R4242 VSS.n4607 VSS.n4606 100.713
R4243 VSS.n4634 VSS.n4607 100.713
R4244 VSS.n4634 VSS.n4633 100.713
R4245 VSS.n4633 VSS.n4632 100.713
R4246 VSS.n4632 VSS.n4608 100.713
R4247 VSS.n4619 VSS.n4618 100.713
R4248 VSS.n4619 VSS.n738 100.713
R4249 VSS.n4646 VSS.n738 100.713
R4250 VSS.n4647 VSS.n4646 100.713
R4251 VSS.n4649 VSS.n4647 100.713
R4252 VSS.n4653 VSS.n565 100.713
R4253 VSS.n5097 VSS.n565 100.713
R4254 VSS.n5097 VSS.n5096 100.713
R4255 VSS.n5096 VSS.n5095 100.713
R4256 VSS.n5095 VSS.n566 100.713
R4257 VSS.n5082 VSS.n574 100.713
R4258 VSS.n5082 VSS.n5081 100.713
R4259 VSS.n5081 VSS.n5080 100.713
R4260 VSS.n5080 VSS.n575 100.713
R4261 VSS.n5070 VSS.n575 100.713
R4262 VSS.n1187 VSS.t72 100.103
R4263 VSS.n5538 VSS.n32 97.5252
R4264 VSS.n4144 VSS.n46 97.5252
R4265 VSS.n5475 VSS.n5474 97.5252
R4266 VSS.n4396 VSS.n1006 97.5252
R4267 VSS.n1523 VSS.n1493 97.5252
R4268 VSS.n2528 VSS.n1558 97.5252
R4269 VSS.n2296 VSS.n2153 97.5252
R4270 VSS.n4654 VSS.n4651 97.5252
R4271 VSS.n4426 VSS.n897 97.5252
R4272 VSS.n4605 VSS.n784 97.5252
R4273 VSS.n3757 VSS.n3583 97.5252
R4274 VSS.n3957 VSS.n1244 97.5252
R4275 VSS.n4019 VSS.n1125 97.5252
R4276 VSS.n5565 VSS.n5564 95.1447
R4277 VSS.n5231 VSS.n5230 93.6243
R4278 VSS.n4951 VSS.n4950 93.6243
R4279 VSS.n610 VSS.n503 93.6243
R4280 VSS.n5040 VSS.n596 93.6243
R4281 VSS.n5257 VSS.n362 93.6243
R4282 VSS.n1219 VSS.n1200 91.7604
R4283 VSS.n1181 VSS.n1170 90.7527
R4284 VSS.n4328 VSS.n1006 89.7233
R4285 VSS.n1493 VSS.n337 89.7233
R4286 VSS.n2535 VSS.n1558 89.7233
R4287 VSS.n2289 VSS.n2153 89.7233
R4288 VSS.n4502 VSS.n784 89.7233
R4289 VSS.n4651 VSS.n4650 89.7233
R4290 VSS.n1244 VSS.n1242 89.7233
R4291 VSS.n1294 VSS.n897 89.7233
R4292 VSS.t62 VSS.t10 87.9115
R4293 VSS.n2994 VSS.n2991 87.7728
R4294 VSS.n3036 VSS.n2991 87.7728
R4295 VSS.n3036 VSS.n2992 87.7728
R4296 VSS.n3032 VSS.n2992 87.7728
R4297 VSS.n3032 VSS.n2997 87.7728
R4298 VSS.n3003 VSS.n2997 87.7728
R4299 VSS.n3003 VSS.n1462 87.7728
R4300 VSS.n3050 VSS.n1462 87.7728
R4301 VSS.n3050 VSS.n1459 87.7728
R4302 VSS.n3054 VSS.n1459 87.7728
R4303 VSS.n2815 VSS.n2813 87.7728
R4304 VSS.n2843 VSS.n2813 87.7728
R4305 VSS.n2843 VSS.n2814 87.7728
R4306 VSS.n2839 VSS.n2814 87.7728
R4307 VSS.n2839 VSS.n1428 87.7728
R4308 VSS.n3112 VSS.n1428 87.7728
R4309 VSS.n3112 VSS.n1425 87.7728
R4310 VSS.n3118 VSS.n1425 87.7728
R4311 VSS.n3118 VSS.n1426 87.7728
R4312 VSS.n1426 VSS.n420 87.7728
R4313 VSS.n3218 VSS.n3217 87.7728
R4314 VSS.n686 VSS.n675 87.7728
R4315 VSS.n2927 VSS.n2591 87.7728
R4316 VSS.n2962 VSS.n2591 87.7728
R4317 VSS.n2962 VSS.n2592 87.7728
R4318 VSS.n2958 VSS.n2592 87.7728
R4319 VSS.n2958 VSS.n2931 87.7728
R4320 VSS.n2931 VSS.n1446 87.7728
R4321 VSS.n3079 VSS.n1446 87.7728
R4322 VSS.n3079 VSS.n1444 87.7728
R4323 VSS.n3084 VSS.n1444 87.7728
R4324 VSS.n3084 VSS.n404 87.7728
R4325 VSS.n943 VSS.n902 87.7728
R4326 VSS.n943 VSS.n942 87.7728
R4327 VSS.n942 VSS.n904 87.7728
R4328 VSS.n914 VSS.n904 87.7728
R4329 VSS.n931 VSS.n914 87.7728
R4330 VSS.n931 VSS.n928 87.7728
R4331 VSS.n928 VSS.n843 87.7728
R4332 VSS.n4545 VSS.n843 87.7728
R4333 VSS.n4545 VSS.n841 87.7728
R4334 VSS.n4549 VSS.n841 87.7728
R4335 VSS.n3709 VSS.n3588 87.7728
R4336 VSS.n1 VSS.t63 87.478
R4337 VSS.n21 VSS.t67 87.1015
R4338 VSS.n1173 VSS.n1172 86.2123
R4339 VSS.n1181 VSS.n1180 83.577
R4340 VSS.n1167 VSS 82.9476
R4341 VSS.n1179 VSS.n1173 82.6783
R4342 VSS.n2293 VSS.n2153 79.9708
R4343 VSS.n1493 VSS.n251 79.9708
R4344 VSS.n2530 VSS.n1558 79.9708
R4345 VSS.n4399 VSS.n1006 79.9708
R4346 VSS.n19 VSS.n18 78.778
R4347 VSS.n17 VSS.n16 78.778
R4348 VSS.n5561 VSS.n5560 76.3222
R4349 VSS.n5534 VSS.n33 76.3222
R4350 VSS.n1136 VSS.n1135 76.3222
R4351 VSS.n5279 VSS.n5278 76.3222
R4352 VSS.n5280 VSS.n5279 76.3222
R4353 VSS.n4992 VSS.n4991 76.3222
R4354 VSS.n5066 VSS.n584 76.3222
R4355 VSS.n611 VSS.n606 76.3222
R4356 VSS.n5255 VSS.n5254 76.3222
R4357 VSS.n614 VSS.n611 76.3222
R4358 VSS.n5067 VSS.n5066 76.3222
R4359 VSS.n1210 VSS.n1209 76.3222
R4360 VSS.n1213 VSS.n1212 76.3222
R4361 VSS.n3995 VSS.n3994 76.3222
R4362 VSS.n1214 VSS.n1202 76.3222
R4363 VSS.n1212 VSS.n1204 76.3222
R4364 VSS.n1210 VSS.n1205 76.3222
R4365 VSS.n4991 VSS.n627 76.3222
R4366 VSS.n5255 VSS.n365 76.3222
R4367 VSS.n1135 VSS.n74 76.3222
R4368 VSS.n5537 VSS.n33 76.3222
R4369 VSS.n5562 VSS.n5561 76.3222
R4370 VSS.n4313 VSS.n4312 76.062
R4371 VSS.n4313 VSS.n4164 76.062
R4372 VSS.n5461 VSS.n5460 76.062
R4373 VSS.n5461 VSS.n110 76.062
R4374 VSS.n4766 VSS.n542 76.062
R4375 VSS.n4706 VSS.n542 76.062
R4376 VSS.n4875 VSS.n519 76.062
R4377 VSS.n4709 VSS.n519 76.062
R4378 VSS.n4561 VSS.n746 76.062
R4379 VSS.n759 VSS.n746 76.062
R4380 VSS.n872 VSS.n871 76.062
R4381 VSS.n4448 VSS.n871 76.062
R4382 VSS.n2059 VSS.n640 76.062
R4383 VSS.n2390 VSS.n640 76.062
R4384 VSS.n2334 VSS.n2333 76.062
R4385 VSS.n2335 VSS.n2334 76.062
R4386 VSS.n2282 VSS.n2281 76.062
R4387 VSS.n2281 VSS.n2280 76.062
R4388 VSS.n2540 VSS.n1467 76.062
R4389 VSS.n1555 VSS.n1467 76.062
R4390 VSS.n5296 VSS.n5295 76.062
R4391 VSS.n5297 VSS.n5296 76.062
R4392 VSS.n4320 VSS.n1019 76.062
R4393 VSS.n4321 VSS.n4320 76.062
R4394 VSS.n1976 VSS.n1975 76.062
R4395 VSS.n1975 VSS.n1974 76.062
R4396 VSS.n3088 VSS.n3087 76.062
R4397 VSS.n3089 VSS.n3088 76.062
R4398 VSS.n2644 VSS.n172 76.062
R4399 VSS.n2637 VSS.n172 76.062
R4400 VSS.n3155 VSS.n849 76.062
R4401 VSS.n1403 VSS.n849 76.062
R4402 VSS.n3842 VSS.n3841 76.062
R4403 VSS.n3843 VSS.n3842 76.062
R4404 VSS.n4061 VSS.n1060 74.5978
R4405 VSS.n3785 VSS.n3784 74.5978
R4406 VSS.n3785 VSS.n3777 74.5978
R4407 VSS.n3648 VSS.n3639 74.5978
R4408 VSS.n3639 VSS.n3638 74.5978
R4409 VSS.n3476 VSS.n3445 74.5978
R4410 VSS.n3445 VSS.n3444 74.5978
R4411 VSS.n4935 VSS.n4821 74.5978
R4412 VSS.n4821 VSS.n4820 74.5978
R4413 VSS.n5176 VSS.n5175 74.5978
R4414 VSS.n5175 VSS.n5174 74.5978
R4415 VSS.n5155 VSS.n449 74.5978
R4416 VSS.n3175 VSS.n449 74.5978
R4417 VSS.n2449 VSS.n2448 74.5978
R4418 VSS.n2448 VSS.n2447 74.5978
R4419 VSS.n2498 VSS.n1579 74.5978
R4420 VSS.n1726 VSS.n1579 74.5978
R4421 VSS.n3040 VSS.n2987 74.5978
R4422 VSS.n2987 VSS.n2986 74.5978
R4423 VSS.n5347 VSS.n5346 74.5978
R4424 VSS.n5346 VSS.n5345 74.5978
R4425 VSS.n2847 VSS.n2809 74.5978
R4426 VSS.n2809 VSS.n2808 74.5978
R4427 VSS.n5409 VSS.n193 74.5978
R4428 VSS.n3351 VSS.n193 74.5978
R4429 VSS.n4062 VSS.n4061 74.5978
R4430 VSS.n5536 VSS.n31 74.0015
R4431 VSS.n1134 VSS.n73 74.0015
R4432 VSS.n3753 VSS.n3752 74.0015
R4433 VSS.n2467 VSS.n1998 73.1441
R4434 VSS.n2175 VSS.n389 73.1441
R4435 VSS.n1918 VSS.n1882 73.1441
R4436 VSS.n1890 VSS.n499 73.1441
R4437 VSS.n4683 VSS.n673 73.1441
R4438 VSS.n291 VSS.n248 73.1441
R4439 VSS.n2593 VSS.n285 73.1441
R4440 VSS.n5374 VSS.n243 73.1441
R4441 VSS.n1346 VSS.n279 73.1441
R4442 VSS.n950 VSS.n266 73.1441
R4443 VSS.n1614 VSS.n1460 73.1441
R4444 VSS.n1623 VSS.n400 73.1441
R4445 VSS.n5191 VSS.n417 73.1441
R4446 VSS.n1388 VSS.n1387 73.1441
R4447 VSS.n3188 VSS.n837 73.1441
R4448 VSS.n1005 VSS.n302 73.1441
R4449 VSS.n4225 VSS.n152 73.1441
R4450 VSS.n3341 VSS.n1004 73.1441
R4451 VSS.n3281 VSS.n3261 73.1441
R4452 VSS.n1003 VSS.n956 73.1441
R4453 VSS.n2995 VSS.n2993 72.8181
R4454 VSS.n2816 VSS.n242 72.8181
R4455 VSS.n2928 VSS.n2926 72.8181
R4456 VSS.n946 VSS.n945 72.8181
R4457 VSS.n1187 VSS.n379 70.5279
R4458 VSS VSS.n5567 70.0568
R4459 VSS.n5565 VSS.n3 67.8811
R4460 VSS.n22 VSS.t92 66.9131
R4461 VSS.n4008 VSS.t89 66.7742
R4462 VSS.n5268 VSS.t72 65.9777
R4463 VSS.t72 VSS.n5244 65.9777
R4464 VSS.n4977 VSS.t72 65.9777
R4465 VSS.n5002 VSS.t72 65.9777
R4466 VSS.n5028 VSS.t72 65.9777
R4467 VSS.n5057 VSS.t72 65.9777
R4468 VSS.t85 VSS.n1049 65.8183
R4469 VSS.t85 VSS.n1047 65.8183
R4470 VSS.t85 VSS.n1045 65.8183
R4471 VSS.n141 VSS.t80 65.8183
R4472 VSS.n5441 VSS.t80 65.8183
R4473 VSS.n5435 VSS.t80 65.8183
R4474 VSS.n5433 VSS.t80 65.8183
R4475 VSS.t74 VSS.n99 65.8183
R4476 VSS.t74 VSS.n97 65.8183
R4477 VSS.t74 VSS.n95 65.8183
R4478 VSS.t53 VSS.n3540 65.8183
R4479 VSS.t53 VSS.n3542 65.8183
R4480 VSS.t53 VSS.n3544 65.8183
R4481 VSS.t53 VSS.n3546 65.8183
R4482 VSS.t53 VSS.n3541 65.8183
R4483 VSS.t53 VSS.n3545 65.8183
R4484 VSS.t53 VSS.n3547 65.8183
R4485 VSS.n3621 VSS.t55 65.8183
R4486 VSS.n3631 VSS.t55 65.8183
R4487 VSS.n3619 VSS.t55 65.8183
R4488 VSS.n3688 VSS.t55 65.8183
R4489 VSS.n3694 VSS.t55 65.8183
R4490 VSS.n3687 VSS.t55 65.8183
R4491 VSS.n3701 VSS.t55 65.8183
R4492 VSS.n3429 VSS.t81 65.8183
R4493 VSS.n3436 VSS.t81 65.8183
R4494 VSS.n3439 VSS.t81 65.8183
R4495 VSS.n3890 VSS.t81 65.8183
R4496 VSS.n1300 VSS.t81 65.8183
R4497 VSS.n3883 VSS.t81 65.8183
R4498 VSS.n3877 VSS.t81 65.8183
R4499 VSS.t73 VSS.n554 65.8183
R4500 VSS.t73 VSS.n552 65.8183
R4501 VSS.t73 VSS.n550 65.8183
R4502 VSS.t73 VSS.n547 65.8183
R4503 VSS.t73 VSS.n551 65.8183
R4504 VSS.t73 VSS.n549 65.8183
R4505 VSS.t73 VSS.n546 65.8183
R4506 VSS.t76 VSS.n531 65.8183
R4507 VSS.t76 VSS.n529 65.8183
R4508 VSS.t76 VSS.n527 65.8183
R4509 VSS.t76 VSS.n524 65.8183
R4510 VSS.t76 VSS.n528 65.8183
R4511 VSS.t76 VSS.n526 65.8183
R4512 VSS.t76 VSS.n523 65.8183
R4513 VSS.n4804 VSS.t79 65.8183
R4514 VSS.n4812 VSS.t79 65.8183
R4515 VSS.n4815 VSS.t79 65.8183
R4516 VSS.n4884 VSS.t79 65.8183
R4517 VSS.n4837 VSS.t79 65.8183
R4518 VSS.n4891 VSS.t79 65.8183
R4519 VSS.n4834 VSS.t79 65.8183
R4520 VSS.n1848 VSS.t75 65.8183
R4521 VSS.n1856 VSS.t75 65.8183
R4522 VSS.n1846 VSS.t75 65.8183
R4523 VSS.n1863 VSS.t75 65.8183
R4524 VSS.n5162 VSS.t75 65.8183
R4525 VSS.n5168 VSS.t75 65.8183
R4526 VSS.n442 VSS.t75 65.8183
R4527 VSS.t58 VSS.n475 65.8183
R4528 VSS.t58 VSS.n477 65.8183
R4529 VSS.t58 VSS.n479 65.8183
R4530 VSS.t58 VSS.n481 65.8183
R4531 VSS.n4640 VSS.t56 65.8183
R4532 VSS.t56 VSS.n772 65.8183
R4533 VSS.t56 VSS.n755 65.8183
R4534 VSS.t56 VSS.n752 65.8183
R4535 VSS.t56 VSS.n756 65.8183
R4536 VSS.t56 VSS.n754 65.8183
R4537 VSS.t56 VSS.n751 65.8183
R4538 VSS.t58 VSS.n476 65.8183
R4539 VSS.t58 VSS.n480 65.8183
R4540 VSS.t58 VSS.n482 65.8183
R4541 VSS.t86 VSS.n885 65.8183
R4542 VSS.t86 VSS.n883 65.8183
R4543 VSS.t86 VSS.n881 65.8183
R4544 VSS.t86 VSS.n878 65.8183
R4545 VSS.t86 VSS.n882 65.8183
R4546 VSS.t86 VSS.n880 65.8183
R4547 VSS.t86 VSS.n877 65.8183
R4548 VSS.n2062 VSS.t99 65.8183
R4549 VSS.n2373 VSS.t99 65.8183
R4550 VSS.n2367 VSS.t99 65.8183
R4551 VSS.n2365 VSS.t99 65.8183
R4552 VSS.n4940 VSS.t96 65.8183
R4553 VSS.t96 VSS.n651 65.8183
R4554 VSS.t96 VSS.n649 65.8183
R4555 VSS.t96 VSS.n646 65.8183
R4556 VSS.t96 VSS.n650 65.8183
R4557 VSS.t96 VSS.n648 65.8183
R4558 VSS.t96 VSS.n645 65.8183
R4559 VSS.n2436 VSS.t99 65.8183
R4560 VSS.n2439 VSS.t99 65.8183
R4561 VSS.n2445 VSS.t99 65.8183
R4562 VSS.n2350 VSS.t71 65.8183
R4563 VSS.n2344 VSS.t71 65.8183
R4564 VSS.n2342 VSS.t71 65.8183
R4565 VSS.n2336 VSS.t71 65.8183
R4566 VSS.n2141 VSS.t71 65.8183
R4567 VSS.n2133 VSS.t71 65.8183
R4568 VSS.n2148 VSS.t71 65.8183
R4569 VSS.n2265 VSS.t98 65.8183
R4570 VSS.n2267 VSS.t98 65.8183
R4571 VSS.n2273 VSS.t98 65.8183
R4572 VSS.n2275 VSS.t98 65.8183
R4573 VSS.n2508 VSS.t98 65.8183
R4574 VSS.n1572 VSS.t98 65.8183
R4575 VSS.n1570 VSS.t98 65.8183
R4576 VSS.n3045 VSS.t84 65.8183
R4577 VSS.t84 VSS.n1478 65.8183
R4578 VSS.t84 VSS.n1476 65.8183
R4579 VSS.t84 VSS.n1473 65.8183
R4580 VSS.t84 VSS.n1477 65.8183
R4581 VSS.t84 VSS.n1475 65.8183
R4582 VSS.t84 VSS.n1472 65.8183
R4583 VSS.n5312 VSS.t78 65.8183
R4584 VSS.n5306 VSS.t78 65.8183
R4585 VSS.n5304 VSS.t78 65.8183
R4586 VSS.n5298 VSS.t78 65.8183
R4587 VSS.n4376 VSS.t78 65.8183
R4588 VSS.n4369 VSS.t78 65.8183
R4589 VSS.n4367 VSS.t78 65.8183
R4590 VSS.t97 VSS.n1032 65.8183
R4591 VSS.t97 VSS.n1030 65.8183
R4592 VSS.t97 VSS.n1028 65.8183
R4593 VSS.t97 VSS.n1025 65.8183
R4594 VSS.n2303 VSS.t71 65.8183
R4595 VSS.n2305 VSS.t71 65.8183
R4596 VSS.n2319 VSS.t71 65.8183
R4597 VSS.n2321 VSS.t71 65.8183
R4598 VSS.n2520 VSS.t98 65.8183
R4599 VSS.n2238 VSS.t98 65.8183
R4600 VSS.n2240 VSS.t98 65.8183
R4601 VSS.n2252 VSS.t98 65.8183
R4602 VSS.t84 VSS.n1471 65.8183
R4603 VSS.t84 VSS.n1470 65.8183
R4604 VSS.t84 VSS.n1469 65.8183
R4605 VSS.t84 VSS.n1468 65.8183
R4606 VSS.n4388 VSS.t78 65.8183
R4607 VSS.n4339 VSS.t78 65.8183
R4608 VSS.n4356 VSS.t78 65.8183
R4609 VSS.n4344 VSS.t78 65.8183
R4610 VSS.t97 VSS.n1021 65.8183
R4611 VSS.t97 VSS.n1022 65.8183
R4612 VSS.t97 VSS.n1023 65.8183
R4613 VSS.t97 VSS.n1024 65.8183
R4614 VSS.t87 VSS.n1599 65.8183
R4615 VSS.t87 VSS.n1601 65.8183
R4616 VSS.t87 VSS.n1603 65.8183
R4617 VSS.t87 VSS.n1605 65.8183
R4618 VSS.n1959 VSS.t83 65.8183
R4619 VSS.n1961 VSS.t83 65.8183
R4620 VSS.n1967 VSS.t83 65.8183
R4621 VSS.n1969 VSS.t83 65.8183
R4622 VSS.n1753 VSS.t83 65.8183
R4623 VSS.n1744 VSS.t83 65.8183
R4624 VSS.n1724 VSS.t83 65.8183
R4625 VSS.t87 VSS.n1600 65.8183
R4626 VSS.t87 VSS.n1604 65.8183
R4627 VSS.t87 VSS.n1606 65.8183
R4628 VSS.n1451 VSS.t77 65.8183
R4629 VSS.n3068 VSS.t77 65.8183
R4630 VSS.n3062 VSS.t77 65.8183
R4631 VSS.n3060 VSS.t77 65.8183
R4632 VSS.n3104 VSS.t68 65.8183
R4633 VSS.n3098 VSS.t68 65.8183
R4634 VSS.n3096 VSS.t68 65.8183
R4635 VSS.n3090 VSS.t68 65.8183
R4636 VSS.n2857 VSS.t68 65.8183
R4637 VSS.n2729 VSS.t68 65.8183
R4638 VSS.n2864 VSS.t68 65.8183
R4639 VSS.n2974 VSS.t77 65.8183
R4640 VSS.n2980 VSS.t77 65.8183
R4641 VSS.n2580 VSS.t77 65.8183
R4642 VSS.n2716 VSS.t70 65.8183
R4643 VSS.n2710 VSS.t70 65.8183
R4644 VSS.n2708 VSS.t70 65.8183
R4645 VSS.n2702 VSS.t70 65.8183
R4646 VSS.t59 VSS.n184 65.8183
R4647 VSS.t59 VSS.n182 65.8183
R4648 VSS.t59 VSS.n180 65.8183
R4649 VSS.t59 VSS.n177 65.8183
R4650 VSS.t59 VSS.n181 65.8183
R4651 VSS.t59 VSS.n179 65.8183
R4652 VSS.t59 VSS.n176 65.8183
R4653 VSS.n5334 VSS.t70 65.8183
R4654 VSS.n5337 VSS.t70 65.8183
R4655 VSS.n5343 VSS.t70 65.8183
R4656 VSS.n2672 VSS.t70 65.8183
R4657 VSS.n2660 VSS.t70 65.8183
R4658 VSS.n2649 VSS.t70 65.8183
R4659 VSS.n5419 VSS.t70 65.8183
R4660 VSS.t59 VSS.n175 65.8183
R4661 VSS.n5414 VSS.t59 65.8183
R4662 VSS.t59 VSS.n174 65.8183
R4663 VSS.t59 VSS.n173 65.8183
R4664 VSS.n3075 VSS.t77 65.8183
R4665 VSS.n2953 VSS.t77 65.8183
R4666 VSS.n2940 VSS.t77 65.8183
R4667 VSS.n2934 VSS.t77 65.8183
R4668 VSS.n2966 VSS.t68 65.8183
R4669 VSS.n2946 VSS.t68 65.8183
R4670 VSS.n2949 VSS.t68 65.8183
R4671 VSS.n2944 VSS.t68 65.8183
R4672 VSS.t87 VSS.n1598 65.8183
R4673 VSS.t87 VSS.n1597 65.8183
R4674 VSS.t87 VSS.n1596 65.8183
R4675 VSS.t87 VSS.n1595 65.8183
R4676 VSS.n1764 VSS.t83 65.8183
R4677 VSS.n1782 VSS.t83 65.8183
R4678 VSS.n1784 VSS.t83 65.8183
R4679 VSS.n1802 VSS.t83 65.8183
R4680 VSS.n2061 VSS.t99 65.8183
R4681 VSS.n2411 VSS.t99 65.8183
R4682 VSS.n2048 VSS.t99 65.8183
R4683 VSS.n2426 VSS.t99 65.8183
R4684 VSS.t96 VSS.n644 65.8183
R4685 VSS.t96 VSS.n643 65.8183
R4686 VSS.t96 VSS.n642 65.8183
R4687 VSS.t96 VSS.n641 65.8183
R4688 VSS.n3139 VSS.t100 65.8183
R4689 VSS.n3133 VSS.t100 65.8183
R4690 VSS.n3131 VSS.t100 65.8183
R4691 VSS.n3125 VSS.t100 65.8183
R4692 VSS.n4540 VSS.t88 65.8183
R4693 VSS.t88 VSS.n860 65.8183
R4694 VSS.t88 VSS.n858 65.8183
R4695 VSS.t88 VSS.n855 65.8183
R4696 VSS.t88 VSS.n859 65.8183
R4697 VSS.t88 VSS.n857 65.8183
R4698 VSS.t88 VSS.n854 65.8183
R4699 VSS.n2796 VSS.t100 65.8183
R4700 VSS.n2802 VSS.t100 65.8183
R4701 VSS.n2739 VSS.t100 65.8183
R4702 VSS.t95 VSS.n209 65.8183
R4703 VSS.t95 VSS.n211 65.8183
R4704 VSS.t95 VSS.n213 65.8183
R4705 VSS.t95 VSS.n215 65.8183
R4706 VSS.n3858 VSS.t82 65.8183
R4707 VSS.n3852 VSS.t82 65.8183
R4708 VSS.n3850 VSS.t82 65.8183
R4709 VSS.n3844 VSS.t82 65.8183
R4710 VSS.n3416 VSS.t82 65.8183
R4711 VSS.n3488 VSS.t82 65.8183
R4712 VSS.n3494 VSS.t82 65.8183
R4713 VSS.t95 VSS.n210 65.8183
R4714 VSS.t95 VSS.n214 65.8183
R4715 VSS.t95 VSS.n216 65.8183
R4716 VSS.t95 VSS.n208 65.8183
R4717 VSS.t95 VSS.n207 65.8183
R4718 VSS.t95 VSS.n206 65.8183
R4719 VSS.t95 VSS.n205 65.8183
R4720 VSS.n3497 VSS.t82 65.8183
R4721 VSS.n3373 VSS.t82 65.8183
R4722 VSS.n3400 VSS.t82 65.8183
R4723 VSS.n3385 VSS.t82 65.8183
R4724 VSS.n3142 VSS.t100 65.8183
R4725 VSS.t100 VSS.n1416 65.8183
R4726 VSS.n2762 VSS.t100 65.8183
R4727 VSS.n2750 VSS.t100 65.8183
R4728 VSS.t88 VSS.n853 65.8183
R4729 VSS.t88 VSS.n852 65.8183
R4730 VSS.t88 VSS.n851 65.8183
R4731 VSS.t88 VSS.n850 65.8183
R4732 VSS.t88 VSS.n846 65.8183
R4733 VSS.t88 VSS.n862 65.8183
R4734 VSS.t88 VSS.n863 65.8183
R4735 VSS.t88 VSS.n864 65.8183
R4736 VSS.n4534 VSS.t86 65.8183
R4737 VSS.t86 VSS.n876 65.8183
R4738 VSS.t86 VSS.n875 65.8183
R4739 VSS.t86 VSS.n874 65.8183
R4740 VSS.t58 VSS.n474 65.8183
R4741 VSS.t58 VSS.n473 65.8183
R4742 VSS.t58 VSS.n472 65.8183
R4743 VSS.t58 VSS.n471 65.8183
R4744 VSS.t56 VSS.n750 65.8183
R4745 VSS.t56 VSS.n749 65.8183
R4746 VSS.t56 VSS.n748 65.8183
R4747 VSS.t56 VSS.n747 65.8183
R4748 VSS.n1849 VSS.t75 65.8183
R4749 VSS.n5142 VSS.t75 65.8183
R4750 VSS.n464 VSS.t75 65.8183
R4751 VSS.n460 VSS.t75 65.8183
R4752 VSS.t58 VSS.n450 65.8183
R4753 VSS.n5133 VSS.t58 65.8183
R4754 VSS.n5137 VSS.t58 65.8183
R4755 VSS.t58 VSS.n5129 65.8183
R4756 VSS.n4853 VSS.t79 65.8183
R4757 VSS.n4856 VSS.t79 65.8183
R4758 VSS.n4844 VSS.t79 65.8183
R4759 VSS.n5114 VSS.t79 65.8183
R4760 VSS.t76 VSS.n522 65.8183
R4761 VSS.n5109 VSS.t76 65.8183
R4762 VSS.t76 VSS.n521 65.8183
R4763 VSS.t76 VSS.n520 65.8183
R4764 VSS.t76 VSS.n532 65.8183
R4765 VSS.t76 VSS.n533 65.8183
R4766 VSS.t76 VSS.n534 65.8183
R4767 VSS.t76 VSS.n535 65.8183
R4768 VSS.n5103 VSS.t73 65.8183
R4769 VSS.t73 VSS.n545 65.8183
R4770 VSS.t73 VSS.n544 65.8183
R4771 VSS.t73 VSS.n543 65.8183
R4772 VSS.t73 VSS.n555 65.8183
R4773 VSS.t73 VSS.n556 65.8183
R4774 VSS.t73 VSS.n557 65.8183
R4775 VSS.t73 VSS.n558 65.8183
R4776 VSS.t56 VSS.n742 65.8183
R4777 VSS.t56 VSS.n774 65.8183
R4778 VSS.t56 VSS.n775 65.8183
R4779 VSS.t56 VSS.n776 65.8183
R4780 VSS.t86 VSS.n886 65.8183
R4781 VSS.t86 VSS.n887 65.8183
R4782 VSS.t86 VSS.n888 65.8183
R4783 VSS.t86 VSS.n889 65.8183
R4784 VSS.n1298 VSS.t81 65.8183
R4785 VSS.n3935 VSS.t81 65.8183
R4786 VSS.n1284 VSS.t81 65.8183
R4787 VSS.n3950 VSS.t81 65.8183
R4788 VSS.n3968 VSS.t55 65.8183
R4789 VSS.n1238 VSS.t55 65.8183
R4790 VSS.n3980 VSS.t55 65.8183
R4791 VSS.t55 VSS.n1225 65.8183
R4792 VSS.t53 VSS.n3539 65.8183
R4793 VSS.t53 VSS.n3538 65.8183
R4794 VSS.t53 VSS.n3537 65.8183
R4795 VSS.t53 VSS.n3536 65.8183
R4796 VSS.n3646 VSS.t55 65.8183
R4797 VSS.n3643 VSS.t55 65.8183
R4798 VSS.n3640 VSS.t55 65.8183
R4799 VSS.n3683 VSS.t55 65.8183
R4800 VSS.n3861 VSS.t82 65.8183
R4801 VSS.t82 VSS.n1317 65.8183
R4802 VSS.n3468 VSS.t82 65.8183
R4803 VSS.n3449 VSS.t82 65.8183
R4804 VSS.n3446 VSS.t81 65.8183
R4805 VSS.n3463 VSS.t81 65.8183
R4806 VSS.n3458 VSS.t81 65.8183
R4807 VSS.n3874 VSS.t81 65.8183
R4808 VSS.t74 VSS.n102 65.8183
R4809 VSS.t74 VSS.n103 65.8183
R4810 VSS.t74 VSS.n104 65.8183
R4811 VSS.t74 VSS.n105 65.8183
R4812 VSS.t53 VSS.n3577 65.8183
R4813 VSS.n3786 VSS.t53 65.8183
R4814 VSS.t53 VSS.n3576 65.8183
R4815 VSS.t53 VSS.n3550 65.8183
R4816 VSS.t74 VSS.n98 65.8183
R4817 VSS.t74 VSS.n96 65.8183
R4818 VSS.t74 VSS.n94 65.8183
R4819 VSS.t74 VSS.n93 65.8183
R4820 VSS.n4050 VSS.t80 65.8183
R4821 VSS.n4053 VSS.t80 65.8183
R4822 VSS.n4059 VSS.t80 65.8183
R4823 VSS.t96 VSS.n637 65.8183
R4824 VSS.t96 VSS.n653 65.8183
R4825 VSS.t96 VSS.n654 65.8183
R4826 VSS.t96 VSS.n655 65.8183
R4827 VSS.n4822 VSS.t79 65.8183
R4828 VSS.n4922 VSS.t79 65.8183
R4829 VSS.n4901 VSS.t79 65.8183
R4830 VSS.n4899 VSS.t79 65.8183
R4831 VSS.n1833 VSS.t83 65.8183
R4832 VSS.n1832 VSS.t83 65.8183
R4833 VSS.n1820 VSS.t83 65.8183
R4834 VSS.n5183 VSS.t83 65.8183
R4835 VSS.n5178 VSS.t75 65.8183
R4836 VSS.n1818 VSS.t75 65.8183
R4837 VSS.n1841 VSS.t75 65.8183
R4838 VSS.n1867 VSS.t75 65.8183
R4839 VSS.n3107 VSS.t68 65.8183
R4840 VSS.t68 VSS.n1432 65.8183
R4841 VSS.n2832 VSS.t68 65.8183
R4842 VSS.n2820 VSS.t68 65.8183
R4843 VSS.n2810 VSS.t100 65.8183
R4844 VSS.n2825 VSS.t100 65.8183
R4845 VSS.n2822 VSS.t100 65.8183
R4846 VSS.n3122 VSS.t100 65.8183
R4847 VSS.t59 VSS.n185 65.8183
R4848 VSS.t59 VSS.n186 65.8183
R4849 VSS.t59 VSS.n187 65.8183
R4850 VSS.t59 VSS.n188 65.8183
R4851 VSS.t95 VSS.n194 65.8183
R4852 VSS.n5396 VSS.t95 65.8183
R4853 VSS.t95 VSS.n5395 65.8183
R4854 VSS.t95 VSS.n218 65.8183
R4855 VSS.n5448 VSS.t80 65.8183
R4856 VSS.n119 VSS.t80 65.8183
R4857 VSS.n122 VSS.t80 65.8183
R4858 VSS.n5467 VSS.t80 65.8183
R4859 VSS.t74 VSS.n107 65.8183
R4860 VSS.n5462 VSS.t74 65.8183
R4861 VSS.t74 VSS.n108 65.8183
R4862 VSS.t74 VSS.n109 65.8183
R4863 VSS.t85 VSS.n1052 65.8183
R4864 VSS.t85 VSS.n1053 65.8183
R4865 VSS.t85 VSS.n1054 65.8183
R4866 VSS.t85 VSS.n4159 65.8183
R4867 VSS.n4154 VSS.t80 65.8183
R4868 VSS.n1070 VSS.t80 65.8183
R4869 VSS.n1095 VSS.t80 65.8183
R4870 VSS.n1098 VSS.t80 65.8183
R4871 VSS.t85 VSS.n1048 65.8183
R4872 VSS.t85 VSS.n1046 65.8183
R4873 VSS.t85 VSS.n1044 65.8183
R4874 VSS.t85 VSS.n1043 65.8183
R4875 VSS.t97 VSS.n1029 65.8183
R4876 VSS.t97 VSS.n1027 65.8183
R4877 VSS.t97 VSS.n1020 65.8183
R4878 VSS.n2109 VSS.t71 65.8183
R4879 VSS.n2095 VSS.t71 65.8183
R4880 VSS.n2084 VSS.t71 65.8183
R4881 VSS.n2456 VSS.t71 65.8183
R4882 VSS.n2451 VSS.t99 65.8183
R4883 VSS.n2082 VSS.t99 65.8183
R4884 VSS.n2103 VSS.t99 65.8183
R4885 VSS.n2080 VSS.t99 65.8183
R4886 VSS.n2261 VSS.t98 65.8183
R4887 VSS.n2258 VSS.t98 65.8183
R4888 VSS.n2488 VSS.t98 65.8183
R4889 VSS.n1588 VSS.t98 65.8183
R4890 VSS.t87 VSS.n1580 65.8183
R4891 VSS.n2483 VSS.t87 65.8183
R4892 VSS.t87 VSS.n2480 65.8183
R4893 VSS.t87 VSS.n1608 65.8183
R4894 VSS.t84 VSS.n1465 65.8183
R4895 VSS.t84 VSS.n1480 65.8183
R4896 VSS.t84 VSS.n1481 65.8183
R4897 VSS.t84 VSS.n1482 65.8183
R4898 VSS.n2988 VSS.t77 65.8183
R4899 VSS.n3012 VSS.t77 65.8183
R4900 VSS.n3024 VSS.t77 65.8183
R4901 VSS.n3015 VSS.t77 65.8183
R4902 VSS.n327 VSS.t78 65.8183
R4903 VSS.n2686 VSS.t78 65.8183
R4904 VSS.n2679 VSS.t78 65.8183
R4905 VSS.n5355 VSS.t78 65.8183
R4906 VSS.n5350 VSS.t70 65.8183
R4907 VSS.n313 VSS.t70 65.8183
R4908 VSS.n2696 VSS.t70 65.8183
R4909 VSS.n2699 VSS.t70 65.8183
R4910 VSS.t97 VSS.n1033 65.8183
R4911 VSS.t97 VSS.n1034 65.8183
R4912 VSS.t97 VSS.n1035 65.8183
R4913 VSS.t97 VSS.n1036 65.8183
R4914 VSS.n4314 VSS.t85 65.8183
R4915 VSS.t85 VSS.n4161 65.8183
R4916 VSS.t85 VSS.n4162 65.8183
R4917 VSS.t85 VSS.n4163 65.8183
R4918 VSS.n5329 VSS.t70 64.1729
R4919 VSS.n2971 VSS.t77 64.1729
R4920 VSS.t87 VSS.n1594 64.1729
R4921 VSS.n2035 VSS.t99 64.1729
R4922 VSS.t95 VSS.n204 64.1729
R4923 VSS.n2793 VSS.t100 64.1729
R4924 VSS.t88 VSS.n4539 64.1729
R4925 VSS.t58 VSS.n470 64.1729
R4926 VSS.n5159 VSS.t75 64.1729
R4927 VSS.n4805 VSS.t79 64.1729
R4928 VSS.t76 VSS.n5108 64.1729
R4929 VSS.t73 VSS.n5102 64.1729
R4930 VSS.t56 VSS.n4639 64.1729
R4931 VSS.t86 VSS.n4533 64.1729
R4932 VSS.t81 VSS.n1276 64.1729
R4933 VSS.n3624 VSS.t55 64.1729
R4934 VSS.t53 VSS.n3535 64.1729
R4935 VSS.n3480 VSS.t82 64.1729
R4936 VSS.t74 VSS.n100 64.1729
R4937 VSS.t96 VSS.n4939 64.1729
R4938 VSS.n1747 VSS.t83 64.1729
R4939 VSS.n2851 VSS.t68 64.1729
R4940 VSS.t59 VSS.n5413 64.1729
R4941 VSS.n1112 VSS.t80 64.1729
R4942 VSS.t85 VSS.n1050 64.1729
R4943 VSS.n2135 VSS.t71 64.1729
R4944 VSS.n2502 VSS.t98 64.1729
R4945 VSS.t84 VSS.n3044 64.1729
R4946 VSS.t78 VSS.n308 64.1729
R4947 VSS.t97 VSS.n4319 64.1729
R4948 VSS.n5538 VSS.n5537 62.4163
R4949 VSS.n5475 VSS.n74 62.4163
R4950 VSS.n5500 VSS.n46 62.4163
R4951 VSS.n4963 VSS.n380 62.4163
R4952 VSS.n4954 VSS.n627 62.4163
R4953 VSS.n5043 VSS.n5041 62.4163
R4954 VSS.n615 VSS.n614 62.4163
R4955 VSS.n365 VSS.n363 62.4163
R4956 VSS.n3724 VSS.n1125 62.4163
R4957 VSS.n3754 VSS.n3583 62.4163
R4958 VSS.n3961 VSS.n963 57.0707
R4959 VSS.n3893 VSS.n247 57.0707
R4960 VSS.n4500 VSS.n343 57.0707
R4961 VSS.n4648 VSS.n345 57.0707
R4962 VSS.n4136 VSS.n1050 56.6572
R4963 VSS.n1112 VSS.n86 56.6572
R4964 VSS.n4026 VSS.n100 56.6572
R4965 VSS.n3650 VSS.n3535 56.6572
R4966 VSS.n3763 VSS.n3535 56.6572
R4967 VSS.n3624 VSS.n3623 56.6572
R4968 VSS.n3625 VSS.n3624 56.6572
R4969 VSS.n3952 VSS.n1276 56.6572
R4970 VSS.n3430 VSS.n1276 56.6572
R4971 VSS.n5102 VSS.n5101 56.6572
R4972 VSS.n5102 VSS.n559 56.6572
R4973 VSS.n5108 VSS.n5107 56.6572
R4974 VSS.n5108 VSS.n536 56.6572
R4975 VSS.n4805 VSS.n512 56.6572
R4976 VSS.n4806 VSS.n4805 56.6572
R4977 VSS.n5159 VSS.n5158 56.6572
R4978 VSS.n5160 VSS.n5159 56.6572
R4979 VSS.n788 VSS.n470 56.6572
R4980 VSS.n4639 VSS.n4638 56.6572
R4981 VSS.n4639 VSS.n777 56.6572
R4982 VSS.n3161 VSS.n470 56.6572
R4983 VSS.n4533 VSS.n4532 56.6572
R4984 VSS.n4533 VSS.n890 56.6572
R4985 VSS.n2428 VSS.n2035 56.6572
R4986 VSS.n4939 VSS.n4938 56.6572
R4987 VSS.n4939 VSS.n656 56.6572
R4988 VSS.n2035 VSS.n2017 56.6572
R4989 VSS.n2135 VSS.n2008 56.6572
R4990 VSS.n2136 VSS.n2135 56.6572
R4991 VSS.n2502 VSS.n2501 56.6572
R4992 VSS.n2503 VSS.n2502 56.6572
R4993 VSS.n3044 VSS.n3043 56.6572
R4994 VSS.n3044 VSS.n1483 56.6572
R4995 VSS.n5357 VSS.n308 56.6572
R4996 VSS.n4371 VSS.n308 56.6572
R4997 VSS.n4319 VSS.n4318 56.6572
R4998 VSS.n1768 VSS.n1594 56.6572
R4999 VSS.n1747 VSS.n431 56.6572
R5000 VSS.n1748 VSS.n1747 56.6572
R5001 VSS.n1740 VSS.n1594 56.6572
R5002 VSS.n2971 VSS.n2970 56.6572
R5003 VSS.n2851 VSS.n2850 56.6572
R5004 VSS.n2852 VSS.n2851 56.6572
R5005 VSS.n2972 VSS.n2971 56.6572
R5006 VSS.n5329 VSS.n165 56.6572
R5007 VSS.n5413 VSS.n5412 56.6572
R5008 VSS.n5413 VSS.n189 56.6572
R5009 VSS.n5330 VSS.n5329 56.6572
R5010 VSS.n2793 VSS.n2792 56.6572
R5011 VSS.n4539 VSS.n4538 56.6572
R5012 VSS.n4539 VSS.n865 56.6572
R5013 VSS.n2794 VSS.n2793 56.6572
R5014 VSS.n3502 VSS.n204 56.6572
R5015 VSS.n3480 VSS.n3479 56.6572
R5016 VSS.n3481 VSS.n3480 56.6572
R5017 VSS.n3365 VSS.n204 56.6572
R5018 VSS.n3779 VSS.n100 56.6572
R5019 VSS.n1113 VSS.n1112 56.6572
R5020 VSS.n4139 VSS.n1050 56.6572
R5021 VSS.n4319 VSS.n1037 56.6572
R5022 VSS.n3959 VSS.n963 55.9517
R5023 VSS.n896 VSS.n247 55.9517
R5024 VSS.n783 VSS.n343 55.9517
R5025 VSS.n4652 VSS.n345 55.9517
R5026 VSS.t58 VSS.n449 55.2026
R5027 VSS.n3639 VSS.t55 55.2026
R5028 VSS.n3445 VSS.t81 55.2026
R5029 VSS.t53 VSS.n3785 55.2026
R5030 VSS.n4821 VSS.t79 55.2026
R5031 VSS.n5175 VSS.t75 55.2026
R5032 VSS.n2809 VSS.t100 55.2026
R5033 VSS.t95 VSS.n193 55.2026
R5034 VSS.n4061 VSS.t80 55.2026
R5035 VSS.n2448 VSS.t99 55.2026
R5036 VSS.t87 VSS.n1579 55.2026
R5037 VSS.n2987 VSS.t77 55.2026
R5038 VSS.n5346 VSS.t70 55.2026
R5039 VSS.n5502 VSS.n5501 55.084
R5040 VSS.n4320 VSS.t97 54.4705
R5041 VSS.n2334 VSS.t71 54.4705
R5042 VSS.n2281 VSS.t98 54.4705
R5043 VSS.t84 VSS.n1467 54.4705
R5044 VSS.n5296 VSS.t78 54.4705
R5045 VSS.t59 VSS.n172 54.4705
R5046 VSS.n3088 VSS.t68 54.4705
R5047 VSS.n1975 VSS.t83 54.4705
R5048 VSS.t96 VSS.n640 54.4705
R5049 VSS.n3842 VSS.t82 54.4705
R5050 VSS.t88 VSS.n849 54.4705
R5051 VSS.t86 VSS.n871 54.4705
R5052 VSS.t56 VSS.n746 54.4705
R5053 VSS.t76 VSS.n519 54.4705
R5054 VSS.t73 VSS.n542 54.4705
R5055 VSS.t74 VSS.n5461 54.4705
R5056 VSS.t85 VSS.n4313 54.4705
R5057 VSS.n4315 VSS.n4314 53.3664
R5058 VSS.n4281 VSS.n4161 53.3664
R5059 VSS.n4289 VSS.n4162 53.3664
R5060 VSS.n4297 VSS.n4163 53.3664
R5061 VSS.n1043 VSS.n1041 53.3664
R5062 VSS.n4124 VSS.n1044 53.3664
R5063 VSS.n4128 VSS.n1046 53.3664
R5064 VSS.n4132 VSS.n1048 53.3664
R5065 VSS.n4159 VSS.n4158 53.3664
R5066 VSS.n1085 VSS.n1054 53.3664
R5067 VSS.n1076 VSS.n1053 53.3664
R5068 VSS.n1101 VSS.n1052 53.3664
R5069 VSS.n4177 VSS.n1045 53.3664
R5070 VSS.n4174 VSS.n1047 53.3664
R5071 VSS.n4170 VSS.n1049 53.3664
R5072 VSS.n4167 VSS.n1049 53.3664
R5073 VSS.n4171 VSS.n1047 53.3664
R5074 VSS.n4175 VSS.n1045 53.3664
R5075 VSS.n5467 VSS.n5466 53.3664
R5076 VSS.n132 VSS.n122 53.3664
R5077 VSS.n140 VSS.n119 53.3664
R5078 VSS.n5448 VSS.n5447 53.3664
R5079 VSS.n5434 VSS.n5433 53.3664
R5080 VSS.n5435 VSS.n143 53.3664
R5081 VSS.n5442 VSS.n5441 53.3664
R5082 VSS.n5446 VSS.n141 53.3664
R5083 VSS.n5443 VSS.n141 53.3664
R5084 VSS.n5441 VSS.n5440 53.3664
R5085 VSS.n5436 VSS.n5435 53.3664
R5086 VSS.n5433 VSS.n5432 53.3664
R5087 VSS.n4154 VSS.n4153 53.3664
R5088 VSS.n1070 VSS.n1059 53.3664
R5089 VSS.n1095 VSS.n1094 53.3664
R5090 VSS.n1098 VSS.n1097 53.3664
R5091 VSS.n4059 VSS.n4058 53.3664
R5092 VSS.n4053 VSS.n1109 53.3664
R5093 VSS.n4050 VSS.n4049 53.3664
R5094 VSS.n4041 VSS.n107 53.3664
R5095 VSS.n5463 VSS.n5462 53.3664
R5096 VSS.n129 VSS.n108 53.3664
R5097 VSS.n137 VSS.n109 53.3664
R5098 VSS.n4042 VSS.n93 53.3664
R5099 VSS.n4038 VSS.n94 53.3664
R5100 VSS.n4034 VSS.n96 53.3664
R5101 VSS.n4030 VSS.n98 53.3664
R5102 VSS.n3791 VSS.n105 53.3664
R5103 VSS.n3556 VSS.n104 53.3664
R5104 VSS.n3570 VSS.n103 53.3664
R5105 VSS.n3562 VSS.n102 53.3664
R5106 VSS.n3509 VSS.n95 53.3664
R5107 VSS.n3513 VSS.n97 53.3664
R5108 VSS.n3517 VSS.n99 53.3664
R5109 VSS.n3519 VSS.n99 53.3664
R5110 VSS.n3516 VSS.n97 53.3664
R5111 VSS.n3512 VSS.n95 53.3664
R5112 VSS.n3659 VSS.n3536 53.3664
R5113 VSS.n3668 VSS.n3537 53.3664
R5114 VSS.n3678 VSS.n3538 53.3664
R5115 VSS.n3606 VSS.n3539 53.3664
R5116 VSS.n3594 VSS.n3546 53.3664
R5117 VSS.n3598 VSS.n3544 53.3664
R5118 VSS.n3602 VSS.n3542 53.3664
R5119 VSS.n3607 VSS.n3540 53.3664
R5120 VSS.n3603 VSS.n3540 53.3664
R5121 VSS.n3599 VSS.n3542 53.3664
R5122 VSS.n3595 VSS.n3544 53.3664
R5123 VSS.n3591 VSS.n3546 53.3664
R5124 VSS.n3778 VSS.n3577 53.3664
R5125 VSS.n3787 VSS.n3786 53.3664
R5126 VSS.n3576 VSS.n3575 53.3664
R5127 VSS.n3566 VSS.n3550 53.3664
R5128 VSS.n3773 VSS.n3547 53.3664
R5129 VSS.n3772 VSS.n3545 53.3664
R5130 VSS.n3764 VSS.n3541 53.3664
R5131 VSS.n3766 VSS.n3541 53.3664
R5132 VSS.n3769 VSS.n3545 53.3664
R5133 VSS.n3776 VSS.n3547 53.3664
R5134 VSS.n3647 VSS.n3646 53.3664
R5135 VSS.n3644 VSS.n3643 53.3664
R5136 VSS.n3641 VSS.n3640 53.3664
R5137 VSS.n3683 VSS.n3682 53.3664
R5138 VSS.n3633 VSS.n3619 53.3664
R5139 VSS.n3631 VSS.n3630 53.3664
R5140 VSS.n3626 VSS.n3621 53.3664
R5141 VSS.n3621 VSS.n3620 53.3664
R5142 VSS.n3632 VSS.n3631 53.3664
R5143 VSS.n3619 VSS.n3617 53.3664
R5144 VSS.n3982 VSS.n1225 53.3664
R5145 VSS.n3980 VSS.n3979 53.3664
R5146 VSS.n1239 VSS.n1238 53.3664
R5147 VSS.n3968 VSS.n3967 53.3664
R5148 VSS.n3701 VSS.n3700 53.3664
R5149 VSS.n3696 VSS.n3687 53.3664
R5150 VSS.n3694 VSS.n3693 53.3664
R5151 VSS.n3689 VSS.n3688 53.3664
R5152 VSS.n3688 VSS.n1240 53.3664
R5153 VSS.n3695 VSS.n3694 53.3664
R5154 VSS.n3687 VSS.n3685 53.3664
R5155 VSS.n3702 VSS.n3701 53.3664
R5156 VSS.n3475 VSS.n3446 53.3664
R5157 VSS.n3463 VSS.n3462 53.3664
R5158 VSS.n3459 VSS.n3458 53.3664
R5159 VSS.n3874 VSS.n3873 53.3664
R5160 VSS.n3439 VSS.n3438 53.3664
R5161 VSS.n3436 VSS.n3435 53.3664
R5162 VSS.n3431 VSS.n3429 53.3664
R5163 VSS.n3429 VSS.n3428 53.3664
R5164 VSS.n3437 VSS.n3436 53.3664
R5165 VSS.n3440 VSS.n3439 53.3664
R5166 VSS.n3950 VSS.n3949 53.3664
R5167 VSS.n3937 VSS.n1284 53.3664
R5168 VSS.n3935 VSS.n3934 53.3664
R5169 VSS.n1299 VSS.n1298 53.3664
R5170 VSS.n3877 VSS.n1302 53.3664
R5171 VSS.n3884 VSS.n3883 53.3664
R5172 VSS.n3888 VSS.n1300 53.3664
R5173 VSS.n3890 VSS.n3889 53.3664
R5174 VSS.n3891 VSS.n3890 53.3664
R5175 VSS.n3885 VSS.n1300 53.3664
R5176 VSS.n3883 VSS.n3882 53.3664
R5177 VSS.n3878 VSS.n3877 53.3664
R5178 VSS.n5090 VSS.n558 53.3664
R5179 VSS.n5087 VSS.n557 53.3664
R5180 VSS.n578 VSS.n556 53.3664
R5181 VSS.n5076 VSS.n555 53.3664
R5182 VSS.n4705 VSS.n547 53.3664
R5183 VSS.n4701 VSS.n550 53.3664
R5184 VSS.n4697 VSS.n552 53.3664
R5185 VSS.n4693 VSS.n554 53.3664
R5186 VSS.n5075 VSS.n554 53.3664
R5187 VSS.n4694 VSS.n552 53.3664
R5188 VSS.n4698 VSS.n550 53.3664
R5189 VSS.n4702 VSS.n547 53.3664
R5190 VSS.n5104 VSS.n5103 53.3664
R5191 VSS.n4744 VSS.n545 53.3664
R5192 VSS.n4752 VSS.n544 53.3664
R5193 VSS.n4760 VSS.n543 53.3664
R5194 VSS.n546 VSS.n540 53.3664
R5195 VSS.n724 VSS.n549 53.3664
R5196 VSS.n728 VSS.n551 53.3664
R5197 VSS.n730 VSS.n551 53.3664
R5198 VSS.n727 VSS.n549 53.3664
R5199 VSS.n721 VSS.n546 53.3664
R5200 VSS.n4747 VSS.n535 53.3664
R5201 VSS.n4755 VSS.n534 53.3664
R5202 VSS.n4763 VSS.n533 53.3664
R5203 VSS.n4771 VSS.n532 53.3664
R5204 VSS.n4710 VSS.n524 53.3664
R5205 VSS.n4714 VSS.n527 53.3664
R5206 VSS.n4718 VSS.n529 53.3664
R5207 VSS.n4722 VSS.n531 53.3664
R5208 VSS.n4772 VSS.n531 53.3664
R5209 VSS.n4721 VSS.n529 53.3664
R5210 VSS.n4717 VSS.n527 53.3664
R5211 VSS.n4713 VSS.n524 53.3664
R5212 VSS.n4797 VSS.n522 53.3664
R5213 VSS.n5110 VSS.n5109 53.3664
R5214 VSS.n4842 VSS.n521 53.3664
R5215 VSS.n4866 VSS.n520 53.3664
R5216 VSS.n4798 VSS.n523 53.3664
R5217 VSS.n4792 VSS.n526 53.3664
R5218 VSS.n4789 VSS.n528 53.3664
R5219 VSS.n4786 VSS.n528 53.3664
R5220 VSS.n4790 VSS.n526 53.3664
R5221 VSS.n4795 VSS.n523 53.3664
R5222 VSS.n4934 VSS.n4822 53.3664
R5223 VSS.n4923 VSS.n4922 53.3664
R5224 VSS.n4901 VSS.n4828 53.3664
R5225 VSS.n4900 VSS.n4899 53.3664
R5226 VSS.n4815 VSS.n4814 53.3664
R5227 VSS.n4812 VSS.n4811 53.3664
R5228 VSS.n4807 VSS.n4804 53.3664
R5229 VSS.n4804 VSS.n667 53.3664
R5230 VSS.n4813 VSS.n4812 53.3664
R5231 VSS.n4816 VSS.n4815 53.3664
R5232 VSS.n5114 VSS.n5113 53.3664
R5233 VSS.n4852 VSS.n4844 53.3664
R5234 VSS.n4856 VSS.n4855 53.3664
R5235 VSS.n4853 VSS.n4838 53.3664
R5236 VSS.n4893 VSS.n4834 53.3664
R5237 VSS.n4891 VSS.n4890 53.3664
R5238 VSS.n4886 VSS.n4837 53.3664
R5239 VSS.n4885 VSS.n4884 53.3664
R5240 VSS.n4884 VSS.n4883 53.3664
R5241 VSS.n4837 VSS.n4835 53.3664
R5242 VSS.n4892 VSS.n4891 53.3664
R5243 VSS.n4834 VSS.n4830 53.3664
R5244 VSS.n461 VSS.n460 53.3664
R5245 VSS.n5144 VSS.n464 53.3664
R5246 VSS.n5142 VSS.n5141 53.3664
R5247 VSS.n1850 VSS.n1849 53.3664
R5248 VSS.n1863 VSS.n1862 53.3664
R5249 VSS.n1858 VSS.n1846 53.3664
R5250 VSS.n1856 VSS.n1855 53.3664
R5251 VSS.n1851 VSS.n1848 53.3664
R5252 VSS.n1848 VSS.n1847 53.3664
R5253 VSS.n1857 VSS.n1856 53.3664
R5254 VSS.n1846 VSS.n1844 53.3664
R5255 VSS.n1864 VSS.n1863 53.3664
R5256 VSS.n5178 VSS.n5177 53.3664
R5257 VSS.n1818 VSS.n436 53.3664
R5258 VSS.n1841 VSS.n1840 53.3664
R5259 VSS.n1868 VSS.n1867 53.3664
R5260 VSS.n5170 VSS.n442 53.3664
R5261 VSS.n5169 VSS.n5168 53.3664
R5262 VSS.n5162 VSS.n5161 53.3664
R5263 VSS.n5163 VSS.n5162 53.3664
R5264 VSS.n5168 VSS.n5167 53.3664
R5265 VSS.n442 VSS.n437 53.3664
R5266 VSS.n4579 VSS.n471 53.3664
R5267 VSS.n806 VSS.n472 53.3664
R5268 VSS.n4566 VSS.n473 53.3664
R5269 VSS.n832 VSS.n474 53.3664
R5270 VSS.n819 VSS.n481 53.3664
R5271 VSS.n823 VSS.n479 53.3664
R5272 VSS.n827 VSS.n477 53.3664
R5273 VSS.n831 VSS.n475 53.3664
R5274 VSS.n828 VSS.n475 53.3664
R5275 VSS.n824 VSS.n477 53.3664
R5276 VSS.n820 VSS.n479 53.3664
R5277 VSS.n816 VSS.n481 53.3664
R5278 VSS.n5154 VSS.n450 53.3664
R5279 VSS.n5133 VSS.n5132 53.3664
R5280 VSS.n5137 VSS.n5136 53.3664
R5281 VSS.n5129 VSS.n469 53.3664
R5282 VSS.n3171 VSS.n482 53.3664
R5283 VSS.n3170 VSS.n480 53.3664
R5284 VSS.n3162 VSS.n476 53.3664
R5285 VSS.n4627 VSS.n776 53.3664
R5286 VSS.n4624 VSS.n775 53.3664
R5287 VSS.n4615 VSS.n774 53.3664
R5288 VSS.n4642 VSS.n742 53.3664
R5289 VSS.n760 VSS.n752 53.3664
R5290 VSS.n764 VSS.n755 53.3664
R5291 VSS.n772 VSS.n757 53.3664
R5292 VSS.n4640 VSS.n745 53.3664
R5293 VSS.n4641 VSS.n4640 53.3664
R5294 VSS.n772 VSS.n771 53.3664
R5295 VSS.n766 VSS.n755 53.3664
R5296 VSS.n763 VSS.n752 53.3664
R5297 VSS.n4587 VSS.n750 53.3664
R5298 VSS.n796 VSS.n749 53.3664
R5299 VSS.n4574 VSS.n748 53.3664
R5300 VSS.n811 VSS.n747 53.3664
R5301 VSS.n4588 VSS.n751 53.3664
R5302 VSS.n4593 VSS.n754 53.3664
R5303 VSS.n4597 VSS.n756 53.3664
R5304 VSS.n4599 VSS.n756 53.3664
R5305 VSS.n4596 VSS.n754 53.3664
R5306 VSS.n4590 VSS.n751 53.3664
R5307 VSS.n3164 VSS.n476 53.3664
R5308 VSS.n3167 VSS.n480 53.3664
R5309 VSS.n3174 VSS.n482 53.3664
R5310 VSS.n4521 VSS.n889 53.3664
R5311 VSS.n4518 VSS.n888 53.3664
R5312 VSS.n4441 VSS.n887 53.3664
R5313 VSS.n4507 VSS.n886 53.3664
R5314 VSS.n4449 VSS.n878 53.3664
R5315 VSS.n4453 VSS.n881 53.3664
R5316 VSS.n4457 VSS.n883 53.3664
R5317 VSS.n4461 VSS.n885 53.3664
R5318 VSS.n4506 VSS.n885 53.3664
R5319 VSS.n4460 VSS.n883 53.3664
R5320 VSS.n4456 VSS.n881 53.3664
R5321 VSS.n4452 VSS.n878 53.3664
R5322 VSS.n4535 VSS.n4534 53.3664
R5323 VSS.n907 VSS.n876 53.3664
R5324 VSS.n934 VSS.n875 53.3664
R5325 VSS.n920 VSS.n874 53.3664
R5326 VSS.n877 VSS.n869 53.3664
R5327 VSS.n4414 VSS.n880 53.3664
R5328 VSS.n4418 VSS.n882 53.3664
R5329 VSS.n4420 VSS.n882 53.3664
R5330 VSS.n4417 VSS.n880 53.3664
R5331 VSS.n4411 VSS.n877 53.3664
R5332 VSS.n2426 VSS.n2425 53.3664
R5333 VSS.n2413 VSS.n2048 53.3664
R5334 VSS.n2411 VSS.n2410 53.3664
R5335 VSS.n2398 VSS.n2061 53.3664
R5336 VSS.n2366 VSS.n2365 53.3664
R5337 VSS.n2367 VSS.n2064 53.3664
R5338 VSS.n2374 VSS.n2373 53.3664
R5339 VSS.n2397 VSS.n2062 53.3664
R5340 VSS.n2375 VSS.n2062 53.3664
R5341 VSS.n2373 VSS.n2372 53.3664
R5342 VSS.n2368 VSS.n2367 53.3664
R5343 VSS.n2365 VSS.n2364 53.3664
R5344 VSS.n2451 VSS.n2450 53.3664
R5345 VSS.n2082 VSS.n2012 53.3664
R5346 VSS.n2103 VSS.n2102 53.3664
R5347 VSS.n2081 VSS.n2080 53.3664
R5348 VSS.n2445 VSS.n2444 53.3664
R5349 VSS.n2439 VSS.n2014 53.3664
R5350 VSS.n2436 VSS.n2435 53.3664
R5351 VSS.n4925 VSS.n655 53.3664
R5352 VSS.n4913 VSS.n654 53.3664
R5353 VSS.n4907 VSS.n653 53.3664
R5354 VSS.n4942 VSS.n637 53.3664
R5355 VSS.n2389 VSS.n646 53.3664
R5356 VSS.n2385 VSS.n649 53.3664
R5357 VSS.n2381 VSS.n651 53.3664
R5358 VSS.n4940 VSS.n639 53.3664
R5359 VSS.n4941 VSS.n4940 53.3664
R5360 VSS.n2378 VSS.n651 53.3664
R5361 VSS.n2382 VSS.n649 53.3664
R5362 VSS.n2386 VSS.n646 53.3664
R5363 VSS.n2033 VSS.n644 53.3664
R5364 VSS.n2422 VSS.n643 53.3664
R5365 VSS.n2046 VSS.n642 53.3664
R5366 VSS.n2407 VSS.n641 53.3664
R5367 VSS.n2032 VSS.n645 53.3664
R5368 VSS.n2026 VSS.n648 53.3664
R5369 VSS.n2023 VSS.n650 53.3664
R5370 VSS.n2020 VSS.n650 53.3664
R5371 VSS.n2024 VSS.n648 53.3664
R5372 VSS.n2029 VSS.n645 53.3664
R5373 VSS.n2437 VSS.n2436 53.3664
R5374 VSS.n2440 VSS.n2439 53.3664
R5375 VSS.n2446 VSS.n2445 53.3664
R5376 VSS.n2456 VSS.n2455 53.3664
R5377 VSS.n2094 VSS.n2084 53.3664
R5378 VSS.n2095 VSS.n2077 53.3664
R5379 VSS.n2352 VSS.n2109 53.3664
R5380 VSS.n2337 VSS.n2336 53.3664
R5381 VSS.n2342 VSS.n2341 53.3664
R5382 VSS.n2345 VSS.n2344 53.3664
R5383 VSS.n2350 VSS.n2349 53.3664
R5384 VSS.n2351 VSS.n2350 53.3664
R5385 VSS.n2344 VSS.n2110 53.3664
R5386 VSS.n2343 VSS.n2342 53.3664
R5387 VSS.n2336 VSS.n2112 53.3664
R5388 VSS.n2303 VSS.n2302 53.3664
R5389 VSS.n2306 VSS.n2305 53.3664
R5390 VSS.n2319 VSS.n2318 53.3664
R5391 VSS.n2322 VSS.n2321 53.3664
R5392 VSS.n2148 VSS.n2131 53.3664
R5393 VSS.n2146 VSS.n2133 53.3664
R5394 VSS.n2142 VSS.n2141 53.3664
R5395 VSS.n2141 VSS.n2140 53.3664
R5396 VSS.n2143 VSS.n2133 53.3664
R5397 VSS.n2149 VSS.n2148 53.3664
R5398 VSS.n1589 VSS.n1588 53.3664
R5399 VSS.n2488 VSS.n2487 53.3664
R5400 VSS.n2259 VSS.n2258 53.3664
R5401 VSS.n2263 VSS.n2261 53.3664
R5402 VSS.n2275 VSS.n2254 53.3664
R5403 VSS.n2274 VSS.n2273 53.3664
R5404 VSS.n2267 VSS.n2256 53.3664
R5405 VSS.n2266 VSS.n2265 53.3664
R5406 VSS.n2265 VSS.n2264 53.3664
R5407 VSS.n2268 VSS.n2267 53.3664
R5408 VSS.n2273 VSS.n2272 53.3664
R5409 VSS.n2276 VSS.n2275 53.3664
R5410 VSS.n2520 VSS.n2519 53.3664
R5411 VSS.n2238 VSS.n1569 53.3664
R5412 VSS.n2241 VSS.n2240 53.3664
R5413 VSS.n2252 VSS.n2251 53.3664
R5414 VSS.n2518 VSS.n1570 53.3664
R5415 VSS.n2513 VSS.n1572 53.3664
R5416 VSS.n2509 VSS.n2508 53.3664
R5417 VSS.n2508 VSS.n2507 53.3664
R5418 VSS.n2510 VSS.n1572 53.3664
R5419 VSS.n2515 VSS.n1570 53.3664
R5420 VSS.n3005 VSS.n1482 53.3664
R5421 VSS.n3029 VSS.n1481 53.3664
R5422 VSS.n3018 VSS.n1480 53.3664
R5423 VSS.n3047 VSS.n1465 53.3664
R5424 VSS.n1554 VSS.n1473 53.3664
R5425 VSS.n1550 VSS.n1476 53.3664
R5426 VSS.n1546 VSS.n1478 53.3664
R5427 VSS.n3045 VSS.n1466 53.3664
R5428 VSS.n3046 VSS.n3045 53.3664
R5429 VSS.n1543 VSS.n1478 53.3664
R5430 VSS.n1547 VSS.n1476 53.3664
R5431 VSS.n1551 VSS.n1473 53.3664
R5432 VSS.n2562 VSS.n1471 53.3664
R5433 VSS.n1530 VSS.n1470 53.3664
R5434 VSS.n2551 VSS.n1469 53.3664
R5435 VSS.n1539 VSS.n1468 53.3664
R5436 VSS.n2563 VSS.n1472 53.3664
R5437 VSS.n2568 VSS.n1475 53.3664
R5438 VSS.n2572 VSS.n1477 53.3664
R5439 VSS.n2574 VSS.n1477 53.3664
R5440 VSS.n2571 VSS.n1475 53.3664
R5441 VSS.n2565 VSS.n1472 53.3664
R5442 VSS.n5355 VSS.n5354 53.3664
R5443 VSS.n2680 VSS.n2679 53.3664
R5444 VSS.n2690 VSS.n2686 53.3664
R5445 VSS.n5314 VSS.n327 53.3664
R5446 VSS.n5299 VSS.n5298 53.3664
R5447 VSS.n5304 VSS.n5303 53.3664
R5448 VSS.n5307 VSS.n5306 53.3664
R5449 VSS.n5312 VSS.n5311 53.3664
R5450 VSS.n5313 VSS.n5312 53.3664
R5451 VSS.n5306 VSS.n329 53.3664
R5452 VSS.n5305 VSS.n5304 53.3664
R5453 VSS.n5298 VSS.n331 53.3664
R5454 VSS.n4388 VSS.n4387 53.3664
R5455 VSS.n4366 VSS.n4339 53.3664
R5456 VSS.n4357 VSS.n4356 53.3664
R5457 VSS.n4345 VSS.n4344 53.3664
R5458 VSS.n4386 VSS.n4367 53.3664
R5459 VSS.n4381 VSS.n4369 53.3664
R5460 VSS.n4377 VSS.n4376 53.3664
R5461 VSS.n4376 VSS.n4375 53.3664
R5462 VSS.n4378 VSS.n4369 53.3664
R5463 VSS.n4383 VSS.n4367 53.3664
R5464 VSS.n4103 VSS.n1021 53.3664
R5465 VSS.n4076 VSS.n1022 53.3664
R5466 VSS.n4092 VSS.n1023 53.3664
R5467 VSS.n4082 VSS.n1024 53.3664
R5468 VSS.n4104 VSS.n1020 53.3664
R5469 VSS.n4109 VSS.n1027 53.3664
R5470 VSS.n4113 VSS.n1029 53.3664
R5471 VSS.n4284 VSS.n1036 53.3664
R5472 VSS.n4292 VSS.n1035 53.3664
R5473 VSS.n4300 VSS.n1034 53.3664
R5474 VSS.n4196 VSS.n1033 53.3664
R5475 VSS.n4182 VSS.n1025 53.3664
R5476 VSS.n4186 VSS.n1028 53.3664
R5477 VSS.n4190 VSS.n1030 53.3664
R5478 VSS.n4194 VSS.n1032 53.3664
R5479 VSS.n4197 VSS.n1032 53.3664
R5480 VSS.n4193 VSS.n1030 53.3664
R5481 VSS.n4189 VSS.n1028 53.3664
R5482 VSS.n4185 VSS.n1025 53.3664
R5483 VSS.n2304 VSS.n2303 53.3664
R5484 VSS.n2305 VSS.n2123 53.3664
R5485 VSS.n2320 VSS.n2319 53.3664
R5486 VSS.n2321 VSS.n2114 53.3664
R5487 VSS.n2521 VSS.n2520 53.3664
R5488 VSS.n2239 VSS.n2238 53.3664
R5489 VSS.n2240 VSS.n2228 53.3664
R5490 VSS.n2253 VSS.n2252 53.3664
R5491 VSS.n1529 VSS.n1471 53.3664
R5492 VSS.n2552 VSS.n1470 53.3664
R5493 VSS.n1538 VSS.n1469 53.3664
R5494 VSS.n2541 VSS.n1468 53.3664
R5495 VSS.n4389 VSS.n4388 53.3664
R5496 VSS.n4343 VSS.n4339 53.3664
R5497 VSS.n4356 VSS.n4355 53.3664
R5498 VSS.n4344 VSS.n333 53.3664
R5499 VSS.n4075 VSS.n1021 53.3664
R5500 VSS.n4093 VSS.n1022 53.3664
R5501 VSS.n4081 VSS.n1023 53.3664
R5502 VSS.n1024 VSS.n1018 53.3664
R5503 VSS.n1775 VSS.n1595 53.3664
R5504 VSS.n1788 VSS.n1596 53.3664
R5505 VSS.n1709 VSS.n1597 53.3664
R5506 VSS.n1979 VSS.n1598 53.3664
R5507 VSS.n1992 VSS.n1605 53.3664
R5508 VSS.n1988 VSS.n1603 53.3664
R5509 VSS.n1984 VSS.n1601 53.3664
R5510 VSS.n1980 VSS.n1599 53.3664
R5511 VSS.n1983 VSS.n1599 53.3664
R5512 VSS.n1987 VSS.n1601 53.3664
R5513 VSS.n1991 VSS.n1603 53.3664
R5514 VSS.n1994 VSS.n1605 53.3664
R5515 VSS.n2497 VSS.n1580 53.3664
R5516 VSS.n2483 VSS.n2482 53.3664
R5517 VSS.n2480 VSS.n1593 53.3664
R5518 VSS.n1609 VSS.n1608 53.3664
R5519 VSS.n1730 VSS.n1606 53.3664
R5520 VSS.n1731 VSS.n1604 53.3664
R5521 VSS.n1739 VSS.n1600 53.3664
R5522 VSS.n5183 VSS.n5182 53.3664
R5523 VSS.n1821 VSS.n1820 53.3664
R5524 VSS.n1835 VSS.n1832 53.3664
R5525 VSS.n1833 VSS.n1808 53.3664
R5526 VSS.n1969 VSS.n1804 53.3664
R5527 VSS.n1968 VSS.n1967 53.3664
R5528 VSS.n1961 VSS.n1806 53.3664
R5529 VSS.n1960 VSS.n1959 53.3664
R5530 VSS.n1959 VSS.n1958 53.3664
R5531 VSS.n1962 VSS.n1961 53.3664
R5532 VSS.n1967 VSS.n1966 53.3664
R5533 VSS.n1970 VSS.n1969 53.3664
R5534 VSS.n1765 VSS.n1764 53.3664
R5535 VSS.n1782 VSS.n1781 53.3664
R5536 VSS.n1785 VSS.n1784 53.3664
R5537 VSS.n1802 VSS.n1801 53.3664
R5538 VSS.n1763 VSS.n1724 53.3664
R5539 VSS.n1758 VSS.n1744 53.3664
R5540 VSS.n1754 VSS.n1753 53.3664
R5541 VSS.n1753 VSS.n1752 53.3664
R5542 VSS.n1755 VSS.n1744 53.3664
R5543 VSS.n1760 VSS.n1724 53.3664
R5544 VSS.n1736 VSS.n1600 53.3664
R5545 VSS.n1733 VSS.n1604 53.3664
R5546 VSS.n1727 VSS.n1606 53.3664
R5547 VSS.n2935 VSS.n2934 53.3664
R5548 VSS.n2955 VSS.n2940 53.3664
R5549 VSS.n2953 VSS.n1450 53.3664
R5550 VSS.n3075 VSS.n3074 53.3664
R5551 VSS.n3061 VSS.n3060 53.3664
R5552 VSS.n3062 VSS.n1453 53.3664
R5553 VSS.n3069 VSS.n3068 53.3664
R5554 VSS.n3073 VSS.n1451 53.3664
R5555 VSS.n3070 VSS.n1451 53.3664
R5556 VSS.n3068 VSS.n3067 53.3664
R5557 VSS.n3063 VSS.n3062 53.3664
R5558 VSS.n3060 VSS.n3059 53.3664
R5559 VSS.n3039 VSS.n2988 53.3664
R5560 VSS.n3012 VSS.n3011 53.3664
R5561 VSS.n3025 VSS.n3024 53.3664
R5562 VSS.n3016 VSS.n3015 53.3664
R5563 VSS.n2982 VSS.n2580 53.3664
R5564 VSS.n2981 VSS.n2980 53.3664
R5565 VSS.n2974 VSS.n2973 53.3664
R5566 VSS.n2821 VSS.n2820 53.3664
R5567 VSS.n2836 VSS.n2832 53.3664
R5568 VSS.n3109 VSS.n1432 53.3664
R5569 VSS.n3107 VSS.n3106 53.3664
R5570 VSS.n3091 VSS.n3090 53.3664
R5571 VSS.n3096 VSS.n3095 53.3664
R5572 VSS.n3099 VSS.n3098 53.3664
R5573 VSS.n3104 VSS.n3103 53.3664
R5574 VSS.n3105 VSS.n3104 53.3664
R5575 VSS.n3098 VSS.n1437 53.3664
R5576 VSS.n3097 VSS.n3096 53.3664
R5577 VSS.n3090 VSS.n1439 53.3664
R5578 VSS.n2967 VSS.n2966 53.3664
R5579 VSS.n2946 VSS.n2588 53.3664
R5580 VSS.n2949 VSS.n2948 53.3664
R5581 VSS.n2945 VSS.n2944 53.3664
R5582 VSS.n2864 VSS.n2587 53.3664
R5583 VSS.n2862 VSS.n2729 53.3664
R5584 VSS.n2858 VSS.n2857 53.3664
R5585 VSS.n2857 VSS.n2856 53.3664
R5586 VSS.n2859 VSS.n2729 53.3664
R5587 VSS.n2865 VSS.n2864 53.3664
R5588 VSS.n2975 VSS.n2974 53.3664
R5589 VSS.n2980 VSS.n2979 53.3664
R5590 VSS.n2580 VSS.n1487 53.3664
R5591 VSS.n5419 VSS.n5418 53.3664
R5592 VSS.n2659 VSS.n2649 53.3664
R5593 VSS.n2660 VSS.n2647 53.3664
R5594 VSS.n2718 VSS.n2672 53.3664
R5595 VSS.n2702 VSS.n2675 53.3664
R5596 VSS.n2709 VSS.n2708 53.3664
R5597 VSS.n2710 VSS.n2673 53.3664
R5598 VSS.n2717 VSS.n2716 53.3664
R5599 VSS.n2716 VSS.n2715 53.3664
R5600 VSS.n2711 VSS.n2710 53.3664
R5601 VSS.n2708 VSS.n2707 53.3664
R5602 VSS.n2703 VSS.n2702 53.3664
R5603 VSS.n5350 VSS.n5349 53.3664
R5604 VSS.n5324 VSS.n313 53.3664
R5605 VSS.n2696 VSS.n2695 53.3664
R5606 VSS.n2699 VSS.n2698 53.3664
R5607 VSS.n5343 VSS.n5342 53.3664
R5608 VSS.n5337 VSS.n5326 53.3664
R5609 VSS.n5334 VSS.n5333 53.3664
R5610 VSS.n5399 VSS.n188 53.3664
R5611 VSS.n225 VSS.n187 53.3664
R5612 VSS.n5385 VSS.n186 53.3664
R5613 VSS.n237 VSS.n185 53.3664
R5614 VSS.n2636 VSS.n177 53.3664
R5615 VSS.n2632 VSS.n180 53.3664
R5616 VSS.n2628 VSS.n182 53.3664
R5617 VSS.n2624 VSS.n184 53.3664
R5618 VSS.n238 VSS.n184 53.3664
R5619 VSS.n2625 VSS.n182 53.3664
R5620 VSS.n2629 VSS.n180 53.3664
R5621 VSS.n2633 VSS.n177 53.3664
R5622 VSS.n3265 VSS.n175 53.3664
R5623 VSS.n5415 VSS.n5414 53.3664
R5624 VSS.n2656 VSS.n174 53.3664
R5625 VSS.n2667 VSS.n173 53.3664
R5626 VSS.n3266 VSS.n176 53.3664
R5627 VSS.n3271 VSS.n179 53.3664
R5628 VSS.n3275 VSS.n181 53.3664
R5629 VSS.n3277 VSS.n181 53.3664
R5630 VSS.n3274 VSS.n179 53.3664
R5631 VSS.n3268 VSS.n176 53.3664
R5632 VSS.n5335 VSS.n5334 53.3664
R5633 VSS.n5338 VSS.n5337 53.3664
R5634 VSS.n5344 VSS.n5343 53.3664
R5635 VSS.n2672 VSS.n2671 53.3664
R5636 VSS.n2661 VSS.n2660 53.3664
R5637 VSS.n2649 VSS.n166 53.3664
R5638 VSS.n5420 VSS.n5419 53.3664
R5639 VSS.n175 VSS.n170 53.3664
R5640 VSS.n5414 VSS.n171 53.3664
R5641 VSS.n2666 VSS.n174 53.3664
R5642 VSS.n2645 VSS.n173 53.3664
R5643 VSS.n3076 VSS.n3075 53.3664
R5644 VSS.n2954 VSS.n2953 53.3664
R5645 VSS.n2940 VSS.n2939 53.3664
R5646 VSS.n2934 VSS.n2584 53.3664
R5647 VSS.n2966 VSS.n2965 53.3664
R5648 VSS.n2947 VSS.n2946 53.3664
R5649 VSS.n2950 VSS.n2949 53.3664
R5650 VSS.n2944 VSS.n1441 53.3664
R5651 VSS.n1710 VSS.n1598 53.3664
R5652 VSS.n1789 VSS.n1597 53.3664
R5653 VSS.n1776 VSS.n1596 53.3664
R5654 VSS.n1769 VSS.n1595 53.3664
R5655 VSS.n1764 VSS.n1719 53.3664
R5656 VSS.n1783 VSS.n1782 53.3664
R5657 VSS.n1784 VSS.n1707 53.3664
R5658 VSS.n1803 VSS.n1802 53.3664
R5659 VSS.n2061 VSS.n2050 53.3664
R5660 VSS.n2412 VSS.n2411 53.3664
R5661 VSS.n2048 VSS.n2037 53.3664
R5662 VSS.n2427 VSS.n2426 53.3664
R5663 VSS.n2421 VSS.n644 53.3664
R5664 VSS.n2045 VSS.n643 53.3664
R5665 VSS.n2406 VSS.n642 53.3664
R5666 VSS.n2058 VSS.n641 53.3664
R5667 VSS.n2751 VSS.n2750 53.3664
R5668 VSS.n2762 VSS.n2761 53.3664
R5669 VSS.n3144 VSS.n1416 53.3664
R5670 VSS.n3142 VSS.n3141 53.3664
R5671 VSS.n3125 VSS.n1419 53.3664
R5672 VSS.n3132 VSS.n3131 53.3664
R5673 VSS.n3133 VSS.n1417 53.3664
R5674 VSS.n3140 VSS.n3139 53.3664
R5675 VSS.n3139 VSS.n3138 53.3664
R5676 VSS.n3134 VSS.n3133 53.3664
R5677 VSS.n3131 VSS.n3130 53.3664
R5678 VSS.n3126 VSS.n3125 53.3664
R5679 VSS.n2846 VSS.n2810 53.3664
R5680 VSS.n2826 VSS.n2825 53.3664
R5681 VSS.n2823 VSS.n2822 53.3664
R5682 VSS.n3122 VSS.n3121 53.3664
R5683 VSS.n2804 VSS.n2739 53.3664
R5684 VSS.n2803 VSS.n2802 53.3664
R5685 VSS.n2796 VSS.n2795 53.3664
R5686 VSS.n939 VSS.n864 53.3664
R5687 VSS.n915 VSS.n863 53.3664
R5688 VSS.n925 VSS.n862 53.3664
R5689 VSS.n4542 VSS.n846 53.3664
R5690 VSS.n1402 VSS.n855 53.3664
R5691 VSS.n1398 VSS.n858 53.3664
R5692 VSS.n1394 VSS.n860 53.3664
R5693 VSS.n4540 VSS.n848 53.3664
R5694 VSS.n4541 VSS.n4540 53.3664
R5695 VSS.n1391 VSS.n860 53.3664
R5696 VSS.n1395 VSS.n858 53.3664
R5697 VSS.n1399 VSS.n855 53.3664
R5698 VSS.n2789 VSS.n853 53.3664
R5699 VSS.n2768 VSS.n852 53.3664
R5700 VSS.n2758 VSS.n851 53.3664
R5701 VSS.n1414 VSS.n850 53.3664
R5702 VSS.n2788 VSS.n854 53.3664
R5703 VSS.n2782 VSS.n857 53.3664
R5704 VSS.n2779 VSS.n859 53.3664
R5705 VSS.n2776 VSS.n859 53.3664
R5706 VSS.n2780 VSS.n857 53.3664
R5707 VSS.n2785 VSS.n854 53.3664
R5708 VSS.n2797 VSS.n2796 53.3664
R5709 VSS.n2802 VSS.n2801 53.3664
R5710 VSS.n2739 VSS.n2737 53.3664
R5711 VSS.n3375 VSS.n205 53.3664
R5712 VSS.n3405 VSS.n206 53.3664
R5713 VSS.n3387 VSS.n207 53.3664
R5714 VSS.n1339 VSS.n208 53.3664
R5715 VSS.n1328 VSS.n215 53.3664
R5716 VSS.n1332 VSS.n213 53.3664
R5717 VSS.n1336 VSS.n211 53.3664
R5718 VSS.n1340 VSS.n209 53.3664
R5719 VSS.n1337 VSS.n209 53.3664
R5720 VSS.n1333 VSS.n211 53.3664
R5721 VSS.n1329 VSS.n213 53.3664
R5722 VSS.n1325 VSS.n215 53.3664
R5723 VSS.n5408 VSS.n194 53.3664
R5724 VSS.n5397 VSS.n5396 53.3664
R5725 VSS.n5395 VSS.n5394 53.3664
R5726 VSS.n5383 VSS.n218 53.3664
R5727 VSS.n3355 VSS.n216 53.3664
R5728 VSS.n3356 VSS.n214 53.3664
R5729 VSS.n3364 VSS.n210 53.3664
R5730 VSS.n3470 VSS.n3449 53.3664
R5731 VSS.n3468 VSS.n3467 53.3664
R5732 VSS.n3863 VSS.n1317 53.3664
R5733 VSS.n3861 VSS.n3860 53.3664
R5734 VSS.n3845 VSS.n3844 53.3664
R5735 VSS.n3850 VSS.n3849 53.3664
R5736 VSS.n3853 VSS.n3852 53.3664
R5737 VSS.n3858 VSS.n3857 53.3664
R5738 VSS.n3859 VSS.n3858 53.3664
R5739 VSS.n3852 VSS.n1319 53.3664
R5740 VSS.n3851 VSS.n3850 53.3664
R5741 VSS.n3844 VSS.n1321 53.3664
R5742 VSS.n3497 VSS.n3496 53.3664
R5743 VSS.n3413 VSS.n3373 53.3664
R5744 VSS.n3400 VSS.n3399 53.3664
R5745 VSS.n3397 VSS.n3385 53.3664
R5746 VSS.n3495 VSS.n3494 53.3664
R5747 VSS.n3489 VSS.n3488 53.3664
R5748 VSS.n3486 VSS.n3416 53.3664
R5749 VSS.n3483 VSS.n3416 53.3664
R5750 VSS.n3488 VSS.n3487 53.3664
R5751 VSS.n3494 VSS.n3493 53.3664
R5752 VSS.n3361 VSS.n210 53.3664
R5753 VSS.n3358 VSS.n214 53.3664
R5754 VSS.n3352 VSS.n216 53.3664
R5755 VSS.n3388 VSS.n208 53.3664
R5756 VSS.n3404 VSS.n207 53.3664
R5757 VSS.n3376 VSS.n206 53.3664
R5758 VSS.n3501 VSS.n205 53.3664
R5759 VSS.n3498 VSS.n3497 53.3664
R5760 VSS.n3398 VSS.n3373 53.3664
R5761 VSS.n3401 VSS.n3400 53.3664
R5762 VSS.n3385 VSS.n1323 53.3664
R5763 VSS.n3143 VSS.n3142 53.3664
R5764 VSS.n2752 VSS.n1416 53.3664
R5765 VSS.n2763 VSS.n2762 53.3664
R5766 VSS.n2750 VSS.n2743 53.3664
R5767 VSS.n2769 VSS.n853 53.3664
R5768 VSS.n2757 VSS.n852 53.3664
R5769 VSS.n1413 VSS.n851 53.3664
R5770 VSS.n3154 VSS.n850 53.3664
R5771 VSS.n924 VSS.n846 53.3664
R5772 VSS.n916 VSS.n862 53.3664
R5773 VSS.n938 VSS.n863 53.3664
R5774 VSS.n866 VSS.n864 53.3664
R5775 VSS.n4534 VSS.n870 53.3664
R5776 VSS.n935 VSS.n876 53.3664
R5777 VSS.n919 VSS.n875 53.3664
R5778 VSS.n874 VSS.n873 53.3664
R5779 VSS.n4565 VSS.n474 53.3664
R5780 VSS.n807 VSS.n473 53.3664
R5781 VSS.n4578 VSS.n472 53.3664
R5782 VSS.n789 VSS.n471 53.3664
R5783 VSS.n795 VSS.n750 53.3664
R5784 VSS.n4575 VSS.n749 53.3664
R5785 VSS.n810 VSS.n748 53.3664
R5786 VSS.n4562 VSS.n747 53.3664
R5787 VSS.n1849 VSS.n466 53.3664
R5788 VSS.n5143 VSS.n5142 53.3664
R5789 VSS.n464 VSS.n463 53.3664
R5790 VSS.n460 VSS.n446 53.3664
R5791 VSS.n5131 VSS.n450 53.3664
R5792 VSS.n5134 VSS.n5133 53.3664
R5793 VSS.n5138 VSS.n5137 53.3664
R5794 VSS.n5129 VSS.n5128 53.3664
R5795 VSS.n4854 VSS.n4853 53.3664
R5796 VSS.n4857 VSS.n4856 53.3664
R5797 VSS.n4844 VSS.n513 53.3664
R5798 VSS.n5115 VSS.n5114 53.3664
R5799 VSS.n522 VSS.n517 53.3664
R5800 VSS.n5109 VSS.n518 53.3664
R5801 VSS.n4865 VSS.n521 53.3664
R5802 VSS.n4874 VSS.n520 53.3664
R5803 VSS.n4764 VSS.n532 53.3664
R5804 VSS.n4756 VSS.n533 53.3664
R5805 VSS.n4748 VSS.n534 53.3664
R5806 VSS.n537 VSS.n535 53.3664
R5807 VSS.n5103 VSS.n541 53.3664
R5808 VSS.n4751 VSS.n545 53.3664
R5809 VSS.n4759 VSS.n544 53.3664
R5810 VSS.n4767 VSS.n543 53.3664
R5811 VSS.n579 VSS.n555 53.3664
R5812 VSS.n5086 VSS.n556 53.3664
R5813 VSS.n5091 VSS.n557 53.3664
R5814 VSS.n560 VSS.n558 53.3664
R5815 VSS.n4614 VSS.n742 53.3664
R5816 VSS.n4623 VSS.n774 53.3664
R5817 VSS.n4628 VSS.n775 53.3664
R5818 VSS.n778 VSS.n776 53.3664
R5819 VSS.n4442 VSS.n886 53.3664
R5820 VSS.n4517 VSS.n887 53.3664
R5821 VSS.n4522 VSS.n888 53.3664
R5822 VSS.n891 VSS.n889 53.3664
R5823 VSS.n1298 VSS.n1286 53.3664
R5824 VSS.n3936 VSS.n3935 53.3664
R5825 VSS.n1284 VSS.n1278 53.3664
R5826 VSS.n3951 VSS.n3950 53.3664
R5827 VSS.n3969 VSS.n3968 53.3664
R5828 VSS.n1238 VSS.n1227 53.3664
R5829 VSS.n3981 VSS.n3980 53.3664
R5830 VSS.n3622 VSS.n1225 53.3664
R5831 VSS.n3679 VSS.n3539 53.3664
R5832 VSS.n3669 VSS.n3538 53.3664
R5833 VSS.n3660 VSS.n3537 53.3664
R5834 VSS.n3651 VSS.n3536 53.3664
R5835 VSS.n3646 VSS.n3645 53.3664
R5836 VSS.n3643 VSS.n3642 53.3664
R5837 VSS.n3640 VSS.n3610 53.3664
R5838 VSS.n3684 VSS.n3683 53.3664
R5839 VSS.n3862 VSS.n3861 53.3664
R5840 VSS.n3453 VSS.n1317 53.3664
R5841 VSS.n3469 VSS.n3468 53.3664
R5842 VSS.n3449 VSS.n3419 53.3664
R5843 VSS.n3460 VSS.n3446 53.3664
R5844 VSS.n3464 VSS.n3463 53.3664
R5845 VSS.n3458 VSS.n1307 53.3664
R5846 VSS.n3875 VSS.n3874 53.3664
R5847 VSS.n3569 VSS.n102 53.3664
R5848 VSS.n3557 VSS.n103 53.3664
R5849 VSS.n3790 VSS.n104 53.3664
R5850 VSS.n3780 VSS.n105 53.3664
R5851 VSS.n3577 VSS.n3533 53.3664
R5852 VSS.n3786 VSS.n3534 53.3664
R5853 VSS.n3576 VSS.n3551 53.3664
R5854 VSS.n3550 VSS.n3549 53.3664
R5855 VSS.n4027 VSS.n98 53.3664
R5856 VSS.n4031 VSS.n96 53.3664
R5857 VSS.n4035 VSS.n94 53.3664
R5858 VSS.n4039 VSS.n93 53.3664
R5859 VSS.n4051 VSS.n4050 53.3664
R5860 VSS.n4054 VSS.n4053 53.3664
R5861 VSS.n4060 VSS.n4059 53.3664
R5862 VSS.n4906 VSS.n637 53.3664
R5863 VSS.n4914 VSS.n653 53.3664
R5864 VSS.n4926 VSS.n654 53.3664
R5865 VSS.n657 VSS.n655 53.3664
R5866 VSS.n4827 VSS.n4822 53.3664
R5867 VSS.n4922 VSS.n4921 53.3664
R5868 VSS.n4902 VSS.n4901 53.3664
R5869 VSS.n4899 VSS.n4898 53.3664
R5870 VSS.n1834 VSS.n1833 53.3664
R5871 VSS.n1832 VSS.n1831 53.3664
R5872 VSS.n1820 VSS.n432 53.3664
R5873 VSS.n5184 VSS.n5183 53.3664
R5874 VSS.n5179 VSS.n5178 53.3664
R5875 VSS.n1819 VSS.n1818 53.3664
R5876 VSS.n1842 VSS.n1841 53.3664
R5877 VSS.n1867 VSS.n1866 53.3664
R5878 VSS.n3108 VSS.n3107 53.3664
R5879 VSS.n2835 VSS.n1432 53.3664
R5880 VSS.n2832 VSS.n2831 53.3664
R5881 VSS.n2820 VSS.n2734 53.3664
R5882 VSS.n2827 VSS.n2810 53.3664
R5883 VSS.n2825 VSS.n2824 53.3664
R5884 VSS.n2822 VSS.n1422 53.3664
R5885 VSS.n3123 VSS.n3122 53.3664
R5886 VSS.n5386 VSS.n185 53.3664
R5887 VSS.n226 VSS.n186 53.3664
R5888 VSS.n5400 VSS.n187 53.3664
R5889 VSS.n190 VSS.n188 53.3664
R5890 VSS.n202 VSS.n194 53.3664
R5891 VSS.n5396 VSS.n203 53.3664
R5892 VSS.n5395 VSS.n219 53.3664
R5893 VSS.n235 VSS.n218 53.3664
R5894 VSS.n5449 VSS.n5448 53.3664
R5895 VSS.n133 VSS.n119 53.3664
R5896 VSS.n122 VSS.n87 53.3664
R5897 VSS.n5468 VSS.n5467 53.3664
R5898 VSS.n107 VSS.n91 53.3664
R5899 VSS.n5462 VSS.n92 53.3664
R5900 VSS.n136 VSS.n108 53.3664
R5901 VSS.n111 VSS.n109 53.3664
R5902 VSS.n1075 VSS.n1052 53.3664
R5903 VSS.n1086 VSS.n1053 53.3664
R5904 VSS.n1056 VSS.n1054 53.3664
R5905 VSS.n4159 VSS.n1055 53.3664
R5906 VSS.n4155 VSS.n4154 53.3664
R5907 VSS.n1071 VSS.n1070 53.3664
R5908 VSS.n1096 VSS.n1095 53.3664
R5909 VSS.n1099 VSS.n1098 53.3664
R5910 VSS.n4135 VSS.n1048 53.3664
R5911 VSS.n4131 VSS.n1046 53.3664
R5912 VSS.n4127 VSS.n1044 53.3664
R5913 VSS.n4123 VSS.n1043 53.3664
R5914 VSS.n4115 VSS.n1029 53.3664
R5915 VSS.n4112 VSS.n1027 53.3664
R5916 VSS.n4106 VSS.n1020 53.3664
R5917 VSS.n2109 VSS.n2108 53.3664
R5918 VSS.n2096 VSS.n2095 53.3664
R5919 VSS.n2084 VSS.n2009 53.3664
R5920 VSS.n2457 VSS.n2456 53.3664
R5921 VSS.n2452 VSS.n2451 53.3664
R5922 VSS.n2083 VSS.n2082 53.3664
R5923 VSS.n2104 VSS.n2103 53.3664
R5924 VSS.n2080 VSS.n2079 53.3664
R5925 VSS.n2261 VSS.n2260 53.3664
R5926 VSS.n2258 VSS.n1590 53.3664
R5927 VSS.n2489 VSS.n2488 53.3664
R5928 VSS.n1588 VSS.n1576 53.3664
R5929 VSS.n2481 VSS.n1580 53.3664
R5930 VSS.n2484 VSS.n2483 53.3664
R5931 VSS.n2480 VSS.n2479 53.3664
R5932 VSS.n1699 VSS.n1608 53.3664
R5933 VSS.n3019 VSS.n1465 53.3664
R5934 VSS.n3028 VSS.n1480 53.3664
R5935 VSS.n3006 VSS.n1481 53.3664
R5936 VSS.n1484 VSS.n1482 53.3664
R5937 VSS.n3010 VSS.n2988 53.3664
R5938 VSS.n3013 VSS.n3012 53.3664
R5939 VSS.n3024 VSS.n3023 53.3664
R5940 VSS.n3015 VSS.n3014 53.3664
R5941 VSS.n2689 VSS.n327 53.3664
R5942 VSS.n2686 VSS.n2685 53.3664
R5943 VSS.n2679 VSS.n310 53.3664
R5944 VSS.n5356 VSS.n5355 53.3664
R5945 VSS.n5351 VSS.n5350 53.3664
R5946 VSS.n2678 VSS.n313 53.3664
R5947 VSS.n2697 VSS.n2696 53.3664
R5948 VSS.n2700 VSS.n2699 53.3664
R5949 VSS.n4301 VSS.n1033 53.3664
R5950 VSS.n4293 VSS.n1034 53.3664
R5951 VSS.n4285 VSS.n1035 53.3664
R5952 VSS.n1038 VSS.n1036 53.3664
R5953 VSS.n4314 VSS.n1042 53.3664
R5954 VSS.n4288 VSS.n4161 53.3664
R5955 VSS.n4296 VSS.n4162 53.3664
R5956 VSS.n4165 VSS.n4163 53.3664
R5957 VSS.n3975 VSS.t54 52.5946
R5958 VSS.n1291 VSS.t60 52.5946
R5959 VSS.n4437 VSS.t69 52.5946
R5960 VSS.n4618 VSS.t57 52.5946
R5961 VSS.t72 VSS.n574 52.5946
R5962 VSS.n5563 VSS.n5 50.0764
R5963 VSS.n5557 VSS.n5556 50.0764
R5964 VSS.n5550 VSS.n5549 50.0764
R5965 VSS.n5549 VSS.n5548 50.0764
R5966 VSS.n5542 VSS.n30 50.0764
R5967 VSS.n5542 VSS.n5541 50.0764
R5968 VSS.n5541 VSS.n5540 50.0764
R5969 VSS.n5536 VSS.n5535 50.0764
R5970 VSS.n5535 VSS.n34 50.0764
R5971 VSS.n38 VSS.n34 50.0764
R5972 VSS.n5528 VSS.n5527 50.0764
R5973 VSS.n5526 VSS.n39 50.0764
R5974 VSS.n5520 VSS.n39 50.0764
R5975 VSS.n5520 VSS.n5519 50.0764
R5976 VSS.n5519 VSS.n5518 50.0764
R5977 VSS.n5518 VSS.n43 50.0764
R5978 VSS.n5512 VSS.n43 50.0764
R5979 VSS.n5495 VSS.n64 50.0764
R5980 VSS.n5494 VSS.n5493 50.0764
R5981 VSS.n5485 VSS.n69 50.0764
R5982 VSS.n5479 VSS.n5478 50.0764
R5983 VSS.n1138 VSS.n1137 50.0764
R5984 VSS.n3726 VSS.n3725 50.0764
R5985 VSS.n3727 VSS.n3726 50.0764
R5986 VSS.n3727 VSS.n3718 50.0764
R5987 VSS.n3733 VSS.n3718 50.0764
R5988 VSS.n3734 VSS.n3733 50.0764
R5989 VSS.n3736 VSS.n3735 50.0764
R5990 VSS.n3744 VSS.n3743 50.0764
R5991 VSS.n3745 VSS.n3744 50.0764
R5992 VSS.n3745 VSS.n3712 50.0764
R5993 VSS.n3751 VSS.n3712 50.0764
R5994 VSS.n3753 VSS.n1192 50.0764
R5995 VSS.n4005 VSS.n1193 50.0764
R5996 VSS.n3999 VSS.n1193 50.0764
R5997 VSS.n3999 VSS.n3998 50.0764
R5998 VSS.n5548 VSS.n26 49.52
R5999 VSS.n5363 VSS.n302 48.7629
R6000 VSS.n2993 VSS.n291 48.7629
R6001 VSS.n5426 VSS.n152 48.7629
R6002 VSS.n3347 VSS.n3341 48.7629
R6003 VSS.n5374 VSS.n242 48.7629
R6004 VSS.n3834 VSS.n3261 48.7629
R6005 VSS.n1682 VSS.n1460 48.7629
R6006 VSS.n5224 VSS.n400 48.7629
R6007 VSS.n5191 VSS.n5190 48.7629
R6008 VSS.n3220 VSS.n1388 48.7629
R6009 VSS.n5228 VSS.n389 48.7629
R6010 VSS.n1918 VSS.n1917 48.7629
R6011 VSS.n5121 VSS.n499 48.7629
R6012 VSS.n4554 VSS.n837 48.7629
R6013 VSS.n4780 VSS.n4683 48.7629
R6014 VSS.n2467 VSS.n2466 48.7629
R6015 VSS.n2926 VSS.n2593 48.7629
R6016 VSS.n3224 VSS.n1346 48.7629
R6017 VSS.n4404 VSS.n956 48.7629
R6018 VSS.n950 VSS.n946 48.7629
R6019 VSS.n1229 VSS.t54 48.1185
R6020 VSS.n3944 VSS.t60 48.1185
R6021 VSS.n4429 VSS.t69 48.1185
R6022 VSS.n4608 VSS.t57 48.1185
R6023 VSS.t72 VSS.n566 48.1185
R6024 VSS.n5558 VSS.t12 47.8508
R6025 VSS.t41 VSS.n1134 47.8508
R6026 VSS.n3735 VSS.t90 47.2944
R6027 VSS.n4006 VSS.n1192 47.2944
R6028 VSS.n4015 VSS.n4014 46.738
R6029 VSS.t44 VSS.n5486 46.1816
R6030 VSS.n5486 VSS.t43 46.1816
R6031 VSS.n710 VSS.t72 45.331
R6032 VSS.n5372 VSS.t69 45.331
R6033 VSS.n407 VSS.t57 45.331
R6034 VSS.n4400 VSS.t60 45.331
R6035 VSS.n4086 VSS.n3 45.1287
R6036 VSS.n4255 VSS.n302 44.8619
R6037 VSS.n152 VSS.n150 44.8619
R6038 VSS.n3341 VSS.n77 44.8619
R6039 VSS.n5365 VSS.n291 44.8619
R6040 VSS.n3054 VSS.n1460 44.8619
R6041 VSS.n2593 VSS.n154 44.8619
R6042 VSS.n5375 VSS.n5374 44.8619
R6043 VSS.n5191 VSS.n420 44.8619
R6044 VSS.n3836 VSS.n1346 44.8619
R6045 VSS.n2468 VSS.n2467 44.8619
R6046 VSS.n5226 VSS.n389 44.8619
R6047 VSS.n1918 VSS.n422 44.8619
R6048 VSS.n5123 VSS.n499 44.8619
R6049 VSS.n4683 VSS.n671 44.8619
R6050 VSS.n404 VSS.n400 44.8619
R6051 VSS.n3222 VSS.n1388 44.8619
R6052 VSS.n4406 VSS.n950 44.8619
R6053 VSS.n4549 VSS.n837 44.8619
R6054 VSS.n960 VSS.n956 44.8619
R6055 VSS.n3261 VSS.n1123 44.8619
R6056 VSS.n674 VSS.t57 44.7423
R6057 VSS.n244 VSS.t60 44.7423
R6058 VSS.n406 VSS.t69 44.7423
R6059 VSS.n1008 VSS.t54 44.7423
R6060 VSS.n55 VSS.t34 42.8976
R6061 VSS.n1164 VSS.t103 42.7603
R6062 VSS.n4010 VSS.t47 42.745
R6063 VSS.n50 VSS.t27 42.6426
R6064 VSS.n1164 VSS.t102 42.6343
R6065 VSS.n50 VSS.t21 42.5516
R6066 VSS.n53 VSS.t24 42.4683
R6067 VSS.n4009 VSS.t46 42.4075
R6068 VSS.n54 VSS.t33 42.3691
R6069 VSS.n5507 VSS.t20 42.3691
R6070 VSS.n5564 VSS.t62 42.2868
R6071 VSS.n25 VSS.n24 41.912
R6072 VSS.n4007 VSS.n4006 41.8265
R6073 VSS.n5540 VSS.n31 41.7304
R6074 VSS.n5477 VSS.n73 41.7304
R6075 VSS.n3722 VSS.n1124 41.7304
R6076 VSS.n3752 VSS.n3751 41.7304
R6077 VSS.n1189 VSS.n1166 41.5908
R6078 VSS.t23 VSS.n1128 41.174
R6079 VSS.n4256 VSS.n32 40.8246
R6080 VSS.n4275 VSS.n4274 40.8246
R6081 VSS.n4274 VSS.n4257 40.8246
R6082 VSS.n4278 VSS.n4277 40.8246
R6083 VSS.n4277 VSS.n4258 40.8246
R6084 VSS.n4272 VSS.n4271 40.8246
R6085 VSS.n4271 VSS.n4259 40.8246
R6086 VSS.n4269 VSS.n4260 40.8246
R6087 VSS.n4306 VSS.n4260 40.8246
R6088 VSS.n4309 VSS.n4200 40.8246
R6089 VSS.n4309 VSS.n4308 40.8246
R6090 VSS.n4144 VSS.n4143 40.8246
R6091 VSS.n4142 VSS.n1062 40.8246
R6092 VSS.n4148 VSS.n4147 40.8246
R6093 VSS.n4147 VSS.n4146 40.8246
R6094 VSS.n1082 VSS.n1081 40.8246
R6095 VSS.n1082 VSS.n1065 40.8246
R6096 VSS.n1091 VSS.n1090 40.8246
R6097 VSS.n1091 VSS.n1066 40.8246
R6098 VSS.n1104 VSS.n1067 40.8246
R6099 VSS.n1107 VSS.n1104 40.8246
R6100 VSS.n1105 VSS.n150 40.8246
R6101 VSS.n5474 VSS.n75 40.8246
R6102 VSS.n5472 VSS.n5471 40.8246
R6103 VSS.n5471 VSS.n83 40.8246
R6104 VSS.n114 VSS.n81 40.8246
R6105 VSS.n115 VSS.n114 40.8246
R6106 VSS.n127 VSS.n80 40.8246
R6107 VSS.n127 VSS.n116 40.8246
R6108 VSS.n117 VSS.n79 40.8246
R6109 VSS.n5454 VSS.n117 40.8246
R6110 VSS.n5457 VSS.n78 40.8246
R6111 VSS.n5457 VSS.n5456 40.8246
R6112 VSS.n5359 VSS.n303 40.8246
R6113 VSS.n318 VSS.n301 40.8246
R6114 VSS.n320 VSS.n319 40.8246
R6115 VSS.n316 VSS.n300 40.8246
R6116 VSS.n5321 VSS.n5320 40.8246
R6117 VSS.n2682 VSS.n299 40.8246
R6118 VSS.n2692 VSS.n321 40.8246
R6119 VSS.n322 VSS.n298 40.8246
R6120 VSS.n5318 VSS.n5317 40.8246
R6121 VSS.n324 VSS.n297 40.8246
R6122 VSS.n5365 VSS.n296 40.8246
R6123 VSS.n159 VSS.n153 40.8246
R6124 VSS.n5424 VSS.n5423 40.8246
R6125 VSS.n167 VSS.n160 40.8246
R6126 VSS.n2640 VSS.n158 40.8246
R6127 VSS.n2652 VSS.n2641 40.8246
R6128 VSS.n2654 VSS.n157 40.8246
R6129 VSS.n2663 VSS.n2642 40.8246
R6130 VSS.n2643 VSS.n156 40.8246
R6131 VSS.n2722 VSS.n2721 40.8246
R6132 VSS.n2725 VSS.n155 40.8246
R6133 VSS.n2724 VSS.n154 40.8246
R6134 VSS.n3346 VSS.n3345 40.8246
R6135 VSS.n3344 VSS.n3343 40.8246
R6136 VSS.n5405 VSS.n197 40.8246
R6137 VSS.n5404 VSS.n5403 40.8246
R6138 VSS.n221 VSS.n199 40.8246
R6139 VSS.n229 VSS.n222 40.8246
R6140 VSS.n5391 VSS.n230 40.8246
R6141 VSS.n5390 VSS.n5389 40.8246
R6142 VSS.n5381 VSS.n231 40.8246
R6143 VSS.n5380 VSS.n5379 40.8246
R6144 VSS.n5375 VSS.n234 40.8246
R6145 VSS.n3504 VSS.n3262 40.8246
R6146 VSS.n3369 VSS.n3260 40.8246
R6147 VSS.n3371 VSS.n3370 40.8246
R6148 VSS.n3410 VSS.n3259 40.8246
R6149 VSS.n3409 VSS.n3408 40.8246
R6150 VSS.n3381 VSS.n3258 40.8246
R6151 VSS.n3383 VSS.n3382 40.8246
R6152 VSS.n3394 VSS.n3257 40.8246
R6153 VSS.n3393 VSS.n3392 40.8246
R6154 VSS.n3838 VSS.n1343 40.8246
R6155 VSS.n3837 VSS.n3836 40.8246
R6156 VSS.n1686 VSS.n1685 40.8246
R6157 VSS.n1684 VSS.n1683 40.8246
R6158 VSS.n2494 VSS.n1583 40.8246
R6159 VSS.n2493 VSS.n2492 40.8246
R6160 VSS.n1687 VSS.n1585 40.8246
R6161 VSS.n1689 VSS.n1688 40.8246
R6162 VSS.n1694 VSS.n1693 40.8246
R6163 VSS.n2476 VSS.n1612 40.8246
R6164 VSS.n2475 VSS.n2474 40.8246
R6165 VSS.n2473 VSS.n2472 40.8246
R6166 VSS.n2468 VSS.n1698 40.8246
R6167 VSS.n1722 VSS.n401 40.8246
R6168 VSS.n1720 VSS.n399 40.8246
R6169 VSS.n1772 VSS.n1712 40.8246
R6170 VSS.n1778 VSS.n398 40.8246
R6171 VSS.n1715 VSS.n1713 40.8246
R6172 VSS.n1714 VSS.n397 40.8246
R6173 VSS.n1794 VSS.n1793 40.8246
R6174 VSS.n1798 VSS.n396 40.8246
R6175 VSS.n1797 VSS.n1796 40.8246
R6176 VSS.n1704 VSS.n395 40.8246
R6177 VSS.n5226 VSS.n394 40.8246
R6178 VSS.n427 VSS.n421 40.8246
R6179 VSS.n5188 VSS.n5187 40.8246
R6180 VSS.n433 VSS.n428 40.8246
R6181 VSS.n1811 VSS.n426 40.8246
R6182 VSS.n1824 VSS.n1812 40.8246
R6183 VSS.n1828 VSS.n425 40.8246
R6184 VSS.n1837 VSS.n1813 40.8246
R6185 VSS.n1814 VSS.n424 40.8246
R6186 VSS.n1873 VSS.n1872 40.8246
R6187 VSS.n1876 VSS.n423 40.8246
R6188 VSS.n1875 VSS.n422 40.8246
R6189 VSS.n3219 VSS.n3218 40.8246
R6190 VSS.n5151 VSS.n453 40.8246
R6191 VSS.n5150 VSS.n5149 40.8246
R6192 VSS.n5148 VSS.n5147 40.8246
R6193 VSS.n487 VSS.n457 40.8246
R6194 VSS.n489 VSS.n488 40.8246
R6195 VSS.n491 VSS.n490 40.8246
R6196 VSS.n496 VSS.n492 40.8246
R6197 VSS.n5125 VSS.n497 40.8246
R6198 VSS.n5125 VSS.n5124 40.8246
R6199 VSS.n2430 VSS.n390 40.8246
R6200 VSS.n2039 VSS.n388 40.8246
R6201 VSS.n2041 VSS.n2040 40.8246
R6202 VSS.n2418 VSS.n387 40.8246
R6203 VSS.n2417 VSS.n2416 40.8246
R6204 VSS.n2052 VSS.n386 40.8246
R6205 VSS.n2054 VSS.n2053 40.8246
R6206 VSS.n2403 VSS.n385 40.8246
R6207 VSS.n2402 VSS.n2401 40.8246
R6208 VSS.n2392 VSS.n384 40.8246
R6209 VSS.n5230 VSS.n382 40.8246
R6210 VSS.n659 VSS.n630 40.8246
R6211 VSS.n661 VSS.n660 40.8246
R6212 VSS.n4931 VSS.n631 40.8246
R6213 VSS.n4930 VSS.n4929 40.8246
R6214 VSS.n4916 VSS.n632 40.8246
R6215 VSS.n4918 VSS.n4917 40.8246
R6216 VSS.n4910 VSS.n633 40.8246
R6217 VSS.n4909 VSS.n634 40.8246
R6218 VSS.n4947 VSS.n4946 40.8246
R6219 VSS.n4945 VSS.n629 40.8246
R6220 VSS.n4950 VSS.n4949 40.8246
R6221 VSS.n508 VSS.n502 40.8246
R6222 VSS.n5119 VSS.n5118 40.8246
R6223 VSS.n514 VSS.n509 40.8246
R6224 VSS.n4847 VSS.n507 40.8246
R6225 VSS.n4849 VSS.n4848 40.8246
R6226 VSS.n4860 VSS.n506 40.8246
R6227 VSS.n4862 VSS.n4861 40.8246
R6228 VSS.n4869 VSS.n505 40.8246
R6229 VSS.n4871 VSS.n4870 40.8246
R6230 VSS.n4879 VSS.n504 40.8246
R6231 VSS.n4878 VSS.n503 40.8246
R6232 VSS.n4553 VSS.n4552 40.8246
R6233 VSS.n4584 VSS.n791 40.8246
R6234 VSS.n4583 VSS.n4582 40.8246
R6235 VSS.n801 VSS.n793 40.8246
R6236 VSS.n803 VSS.n802 40.8246
R6237 VSS.n4571 VSS.n804 40.8246
R6238 VSS.n4570 VSS.n4569 40.8246
R6239 VSS.n834 VSS.n805 40.8246
R6240 VSS.n836 VSS.n835 40.8246
R6241 VSS.n4558 VSS.n4556 40.8246
R6242 VSS.n4558 VSS.n4557 40.8246
R6243 VSS.n4685 VSS.n4684 40.8246
R6244 VSS.n4731 VSS.n4686 40.8246
R6245 VSS.n4742 VSS.n4741 40.8246
R6246 VSS.n4737 VSS.n4687 40.8246
R6247 VSS.n4739 VSS.n4738 40.8246
R6248 VSS.n4734 VSS.n4688 40.8246
R6249 VSS.n4736 VSS.n4735 40.8246
R6250 VSS.n4732 VSS.n4689 40.8246
R6251 VSS.n4733 VSS.n4690 40.8246
R6252 VSS.n4778 VSS.n4777 40.8246
R6253 VSS.n4691 VSS.n596 40.8246
R6254 VSS.n2292 VSS.n2221 40.8246
R6255 VSS.n2220 VSS.n2219 40.8246
R6256 VSS.n2218 VSS.n2217 40.8246
R6257 VSS.n2214 VSS.n2156 40.8246
R6258 VSS.n2213 VSS.n2212 40.8246
R6259 VSS.n2211 VSS.n2210 40.8246
R6260 VSS.n2209 VSS.n2208 40.8246
R6261 VSS.n2205 VSS.n2159 40.8246
R6262 VSS.n2204 VSS.n2203 40.8246
R6263 VSS.n2202 VSS.n2201 40.8246
R6264 VSS.n2201 VSS.n2163 40.8246
R6265 VSS.n2161 VSS.n1998 40.8246
R6266 VSS.n2166 VSS.n2165 40.8246
R6267 VSS.n2197 VSS.n2167 40.8246
R6268 VSS.n2196 VSS.n2195 40.8246
R6269 VSS.n2194 VSS.n2193 40.8246
R6270 VSS.n2192 VSS.n2191 40.8246
R6271 VSS.n2188 VSS.n2169 40.8246
R6272 VSS.n2187 VSS.n2186 40.8246
R6273 VSS.n2185 VSS.n2184 40.8246
R6274 VSS.n2183 VSS.n2182 40.8246
R6275 VSS.n2179 VSS.n2172 40.8246
R6276 VSS.n2179 VSS.n2178 40.8246
R6277 VSS.n2176 VSS.n2175 40.8246
R6278 VSS.n1928 VSS.n1927 40.8246
R6279 VSS.n1930 VSS.n1929 40.8246
R6280 VSS.n1933 VSS.n1924 40.8246
R6281 VSS.n1935 VSS.n1934 40.8246
R6282 VSS.n1937 VSS.n1936 40.8246
R6283 VSS.n1940 VSS.n1922 40.8246
R6284 VSS.n1942 VSS.n1941 40.8246
R6285 VSS.n1944 VSS.n1943 40.8246
R6286 VSS.n1947 VSS.n1920 40.8246
R6287 VSS.n1949 VSS.n1948 40.8246
R6288 VSS.n1950 VSS.n1949 40.8246
R6289 VSS.n1882 VSS.n1878 40.8246
R6290 VSS.n1915 VSS.n1879 40.8246
R6291 VSS.n1914 VSS.n1913 40.8246
R6292 VSS.n1912 VSS.n1911 40.8246
R6293 VSS.n1908 VSS.n1883 40.8246
R6294 VSS.n1907 VSS.n1906 40.8246
R6295 VSS.n1905 VSS.n1904 40.8246
R6296 VSS.n1903 VSS.n1902 40.8246
R6297 VSS.n1899 VSS.n1886 40.8246
R6298 VSS.n1898 VSS.n1897 40.8246
R6299 VSS.n1896 VSS.n1895 40.8246
R6300 VSS.n1895 VSS.n1894 40.8246
R6301 VSS.n1890 VSS.n1889 40.8246
R6302 VSS.n680 VSS.n675 40.8246
R6303 VSS.n689 VSS.n676 40.8246
R6304 VSS.n691 VSS.n690 40.8246
R6305 VSS.n694 VSS.n677 40.8246
R6306 VSS.n696 VSS.n695 40.8246
R6307 VSS.n699 VSS.n678 40.8246
R6308 VSS.n701 VSS.n700 40.8246
R6309 VSS.n703 VSS.n679 40.8246
R6310 VSS.n708 VSS.n684 40.8246
R6311 VSS.n709 VSS.n708 40.8246
R6312 VSS.n682 VSS.n673 40.8246
R6313 VSS.n4681 VSS.n4680 40.8246
R6314 VSS.n4677 VSS.n711 40.8246
R6315 VSS.n4676 VSS.n4675 40.8246
R6316 VSS.n4674 VSS.n4673 40.8246
R6317 VSS.n4672 VSS.n4671 40.8246
R6318 VSS.n4668 VSS.n714 40.8246
R6319 VSS.n4667 VSS.n4666 40.8246
R6320 VSS.n4665 VSS.n4664 40.8246
R6321 VSS.n4663 VSS.n4662 40.8246
R6322 VSS.n4659 VSS.n717 40.8246
R6323 VSS.n4659 VSS.n4658 40.8246
R6324 VSS.n720 VSS.n719 40.8246
R6325 VSS.n4662 VSS.n717 40.8246
R6326 VSS.n4666 VSS.n4665 40.8246
R6327 VSS.n4671 VSS.n714 40.8246
R6328 VSS.n4675 VSS.n4674 40.8246
R6329 VSS.n1897 VSS.n1896 40.8246
R6330 VSS.n1902 VSS.n1886 40.8246
R6331 VSS.n1906 VSS.n1905 40.8246
R6332 VSS.n1911 VSS.n1883 40.8246
R6333 VSS.n1948 VSS.n1947 40.8246
R6334 VSS.n1943 VSS.n1942 40.8246
R6335 VSS.n1937 VSS.n1922 40.8246
R6336 VSS.n1934 VSS.n1933 40.8246
R6337 VSS.n2182 VSS.n2172 40.8246
R6338 VSS.n2186 VSS.n2185 40.8246
R6339 VSS.n2191 VSS.n2169 40.8246
R6340 VSS.n2195 VSS.n2194 40.8246
R6341 VSS.n2203 VSS.n2202 40.8246
R6342 VSS.n2208 VSS.n2159 40.8246
R6343 VSS.n2212 VSS.n2211 40.8246
R6344 VSS.n2217 VSS.n2156 40.8246
R6345 VSS.n2221 VSS.n2220 40.8246
R6346 VSS.n2293 VSS.n2292 40.8246
R6347 VSS.n4664 VSS.n4663 40.8246
R6348 VSS.n4668 VSS.n4667 40.8246
R6349 VSS.n4673 VSS.n4672 40.8246
R6350 VSS.n4677 VSS.n4676 40.8246
R6351 VSS.n1899 VSS.n1898 40.8246
R6352 VSS.n1904 VSS.n1903 40.8246
R6353 VSS.n1908 VSS.n1907 40.8246
R6354 VSS.n1913 VSS.n1912 40.8246
R6355 VSS.n1944 VSS.n1920 40.8246
R6356 VSS.n1941 VSS.n1940 40.8246
R6357 VSS.n1936 VSS.n1935 40.8246
R6358 VSS.n1930 VSS.n1924 40.8246
R6359 VSS.n2184 VSS.n2183 40.8246
R6360 VSS.n2188 VSS.n2187 40.8246
R6361 VSS.n2193 VSS.n2192 40.8246
R6362 VSS.n2197 VSS.n2196 40.8246
R6363 VSS.n2205 VSS.n2204 40.8246
R6364 VSS.n2210 VSS.n2209 40.8246
R6365 VSS.n2214 VSS.n2213 40.8246
R6366 VSS.n2219 VSS.n2218 40.8246
R6367 VSS.n2462 VSS.n2000 40.8246
R6368 VSS.n2461 VSS.n2460 40.8246
R6369 VSS.n2070 VSS.n2005 40.8246
R6370 VSS.n2072 VSS.n2071 40.8246
R6371 VSS.n2088 VSS.n2073 40.8246
R6372 VSS.n2090 VSS.n2089 40.8246
R6373 VSS.n2099 VSS.n2074 40.8246
R6374 VSS.n2098 VSS.n2075 40.8246
R6375 VSS.n2356 VSS.n2355 40.8246
R6376 VSS.n2359 VSS.n2069 40.8246
R6377 VSS.n2358 VSS.n362 40.8246
R6378 VSS.n2392 VSS.n382 40.8246
R6379 VSS.n2401 VSS.n384 40.8246
R6380 VSS.n2403 VSS.n2402 40.8246
R6381 VSS.n2054 VSS.n385 40.8246
R6382 VSS.n2053 VSS.n2052 40.8246
R6383 VSS.n2416 VSS.n386 40.8246
R6384 VSS.n2418 VSS.n2417 40.8246
R6385 VSS.n2041 VSS.n387 40.8246
R6386 VSS.n2040 VSS.n2039 40.8246
R6387 VSS.n2430 VSS.n388 40.8246
R6388 VSS.n1929 VSS.n1928 40.8246
R6389 VSS.n2177 VSS.n2176 40.8246
R6390 VSS.n1927 VSS.n1926 40.8246
R6391 VSS.n2178 VSS.n2177 40.8246
R6392 VSS.n5228 VSS.n390 40.8246
R6393 VSS.n1704 VSS.n394 40.8246
R6394 VSS.n1796 VSS.n395 40.8246
R6395 VSS.n1798 VSS.n1797 40.8246
R6396 VSS.n1793 VSS.n396 40.8246
R6397 VSS.n1794 VSS.n1714 40.8246
R6398 VSS.n1715 VSS.n397 40.8246
R6399 VSS.n1778 VSS.n1713 40.8246
R6400 VSS.n1772 VSS.n398 40.8246
R6401 VSS.n1720 VSS.n1712 40.8246
R6402 VSS.n1722 VSS.n399 40.8246
R6403 VSS.n5224 VSS.n401 40.8246
R6404 VSS.n3224 VSS.n1348 40.8246
R6405 VSS.n2772 VSS.n1349 40.8246
R6406 VSS.n2772 VSS.n1408 40.8246
R6407 VSS.n2765 VSS.n1350 40.8246
R6408 VSS.n2765 VSS.n1409 40.8246
R6409 VSS.n1410 VSS.n1351 40.8246
R6410 VSS.n3148 VSS.n1410 40.8246
R6411 VSS.n1407 VSS.n1352 40.8246
R6412 VSS.n3150 VSS.n1407 40.8246
R6413 VSS.n3157 VSS.n1353 40.8246
R6414 VSS.n3222 VSS.n1354 40.8246
R6415 VSS.n3157 VSS.n1354 40.8246
R6416 VSS.n3151 VSS.n3150 40.8246
R6417 VSS.n3151 VSS.n1353 40.8246
R6418 VSS.n3148 VSS.n3147 40.8246
R6419 VSS.n3147 VSS.n1352 40.8246
R6420 VSS.n2753 VSS.n1409 40.8246
R6421 VSS.n2753 VSS.n1351 40.8246
R6422 VSS.n2746 VSS.n1408 40.8246
R6423 VSS.n2746 VSS.n1350 40.8246
R6424 VSS.n2744 VSS.n1348 40.8246
R6425 VSS.n2744 VSS.n1349 40.8246
R6426 VSS.n4556 VSS.n836 40.8246
R6427 VSS.n835 VSS.n834 40.8246
R6428 VSS.n4569 VSS.n805 40.8246
R6429 VSS.n4571 VSS.n4570 40.8246
R6430 VSS.n804 VSS.n803 40.8246
R6431 VSS.n802 VSS.n801 40.8246
R6432 VSS.n4582 VSS.n793 40.8246
R6433 VSS.n4584 VSS.n4583 40.8246
R6434 VSS.n4552 VSS.n791 40.8246
R6435 VSS.n4554 VSS.n4553 40.8246
R6436 VSS.n3420 VSS.n957 40.8246
R6437 VSS.n3422 VSS.n955 40.8246
R6438 VSS.n3472 VSS.n1311 40.8246
R6439 VSS.n3450 VSS.n954 40.8246
R6440 VSS.n3454 VSS.n1312 40.8246
R6441 VSS.n1313 VSS.n953 40.8246
R6442 VSS.n3867 VSS.n3866 40.8246
R6443 VSS.n1310 VSS.n952 40.8246
R6444 VSS.n3870 VSS.n3869 40.8246
R6445 VSS.n1304 VSS.n951 40.8246
R6446 VSS.n4406 VSS.n948 40.8246
R6447 VSS.n1518 VSS.n290 40.8246
R6448 VSS.n1515 VSS.n1514 40.8246
R6449 VSS.n1512 VSS.n289 40.8246
R6450 VSS.n1511 VSS.n1510 40.8246
R6451 VSS.n1507 VSS.n288 40.8246
R6452 VSS.n1506 VSS.n1505 40.8246
R6453 VSS.n1502 VSS.n287 40.8246
R6454 VSS.n1501 VSS.n1500 40.8246
R6455 VSS.n1497 VSS.n286 40.8246
R6456 VSS.n1496 VSS.n1495 40.8246
R6457 VSS.n1495 VSS.n252 40.8246
R6458 VSS.n5368 VSS.n248 40.8246
R6459 VSS.n292 VSS.n249 40.8246
R6460 VSS.n2595 VSS.n2594 40.8246
R6461 VSS.n2598 VSS.n253 40.8246
R6462 VSS.n2600 VSS.n2599 40.8246
R6463 VSS.n2603 VSS.n254 40.8246
R6464 VSS.n2605 VSS.n2604 40.8246
R6465 VSS.n2608 VSS.n255 40.8246
R6466 VSS.n2610 VSS.n2609 40.8246
R6467 VSS.n2613 VSS.n256 40.8246
R6468 VSS.n2615 VSS.n2614 40.8246
R6469 VSS.n2618 VSS.n257 40.8246
R6470 VSS.n2617 VSS.n285 40.8246
R6471 VSS.n2921 VSS.n284 40.8246
R6472 VSS.n2920 VSS.n2919 40.8246
R6473 VSS.n2916 VSS.n283 40.8246
R6474 VSS.n2915 VSS.n2914 40.8246
R6475 VSS.n2911 VSS.n282 40.8246
R6476 VSS.n2910 VSS.n2909 40.8246
R6477 VSS.n2906 VSS.n281 40.8246
R6478 VSS.n2905 VSS.n2904 40.8246
R6479 VSS.n2901 VSS.n280 40.8246
R6480 VSS.n2900 VSS.n2899 40.8246
R6481 VSS.n2899 VSS.n260 40.8246
R6482 VSS.n258 VSS.n243 40.8246
R6483 VSS.n250 VSS.n245 40.8246
R6484 VSS.n2895 VSS.n2894 40.8246
R6485 VSS.n2892 VSS.n261 40.8246
R6486 VSS.n2891 VSS.n2890 40.8246
R6487 VSS.n2887 VSS.n262 40.8246
R6488 VSS.n2886 VSS.n2885 40.8246
R6489 VSS.n2882 VSS.n263 40.8246
R6490 VSS.n2881 VSS.n2880 40.8246
R6491 VSS.n2877 VSS.n264 40.8246
R6492 VSS.n2876 VSS.n2875 40.8246
R6493 VSS.n2872 VSS.n265 40.8246
R6494 VSS.n2871 VSS.n279 40.8246
R6495 VSS.n3252 VSS.n278 40.8246
R6496 VSS.n3251 VSS.n3250 40.8246
R6497 VSS.n3247 VSS.n277 40.8246
R6498 VSS.n3246 VSS.n3245 40.8246
R6499 VSS.n3242 VSS.n276 40.8246
R6500 VSS.n3241 VSS.n3240 40.8246
R6501 VSS.n3237 VSS.n275 40.8246
R6502 VSS.n3236 VSS.n3235 40.8246
R6503 VSS.n3232 VSS.n274 40.8246
R6504 VSS.n3231 VSS.n3230 40.8246
R6505 VSS.n3227 VSS.n273 40.8246
R6506 VSS.n3226 VSS.n266 40.8246
R6507 VSS.n3898 VSS.n267 40.8246
R6508 VSS.n3900 VSS.n3899 40.8246
R6509 VSS.n3903 VSS.n268 40.8246
R6510 VSS.n3905 VSS.n3904 40.8246
R6511 VSS.n3908 VSS.n269 40.8246
R6512 VSS.n3910 VSS.n3909 40.8246
R6513 VSS.n3913 VSS.n270 40.8246
R6514 VSS.n3915 VSS.n3914 40.8246
R6515 VSS.n3918 VSS.n271 40.8246
R6516 VSS.n3920 VSS.n3919 40.8246
R6517 VSS.n3920 VSS.n272 40.8246
R6518 VSS.n3896 VSS.n3894 40.8246
R6519 VSS.n3919 VSS.n3918 40.8246
R6520 VSS.n3914 VSS.n3913 40.8246
R6521 VSS.n3909 VSS.n3908 40.8246
R6522 VSS.n3904 VSS.n3903 40.8246
R6523 VSS.n3899 VSS.n3898 40.8246
R6524 VSS.n3227 VSS.n3226 40.8246
R6525 VSS.n3232 VSS.n3231 40.8246
R6526 VSS.n3237 VSS.n3236 40.8246
R6527 VSS.n3242 VSS.n3241 40.8246
R6528 VSS.n3247 VSS.n3246 40.8246
R6529 VSS.n3252 VSS.n3251 40.8246
R6530 VSS.n2872 VSS.n2871 40.8246
R6531 VSS.n2877 VSS.n2876 40.8246
R6532 VSS.n2882 VSS.n2881 40.8246
R6533 VSS.n2887 VSS.n2886 40.8246
R6534 VSS.n2892 VSS.n2891 40.8246
R6535 VSS.n2901 VSS.n2900 40.8246
R6536 VSS.n2906 VSS.n2905 40.8246
R6537 VSS.n2911 VSS.n2910 40.8246
R6538 VSS.n2916 VSS.n2915 40.8246
R6539 VSS.n2921 VSS.n2920 40.8246
R6540 VSS.n2618 VSS.n2617 40.8246
R6541 VSS.n2614 VSS.n2613 40.8246
R6542 VSS.n2609 VSS.n2608 40.8246
R6543 VSS.n2604 VSS.n2603 40.8246
R6544 VSS.n2599 VSS.n2598 40.8246
R6545 VSS.n1497 VSS.n1496 40.8246
R6546 VSS.n1502 VSS.n1501 40.8246
R6547 VSS.n1507 VSS.n1506 40.8246
R6548 VSS.n1512 VSS.n1511 40.8246
R6549 VSS.n1514 VSS.n290 40.8246
R6550 VSS.n1518 VSS.n251 40.8246
R6551 VSS.n3915 VSS.n271 40.8246
R6552 VSS.n3910 VSS.n270 40.8246
R6553 VSS.n3905 VSS.n269 40.8246
R6554 VSS.n3900 VSS.n268 40.8246
R6555 VSS.n949 VSS.n267 40.8246
R6556 VSS.n3230 VSS.n273 40.8246
R6557 VSS.n3235 VSS.n274 40.8246
R6558 VSS.n3240 VSS.n275 40.8246
R6559 VSS.n3245 VSS.n276 40.8246
R6560 VSS.n3250 VSS.n277 40.8246
R6561 VSS.n3254 VSS.n278 40.8246
R6562 VSS.n2875 VSS.n265 40.8246
R6563 VSS.n2880 VSS.n264 40.8246
R6564 VSS.n2885 VSS.n263 40.8246
R6565 VSS.n2890 VSS.n262 40.8246
R6566 VSS.n2895 VSS.n261 40.8246
R6567 VSS.n2904 VSS.n280 40.8246
R6568 VSS.n2909 VSS.n281 40.8246
R6569 VSS.n2914 VSS.n282 40.8246
R6570 VSS.n2919 VSS.n283 40.8246
R6571 VSS.n2923 VSS.n284 40.8246
R6572 VSS.n2615 VSS.n257 40.8246
R6573 VSS.n2610 VSS.n256 40.8246
R6574 VSS.n2605 VSS.n255 40.8246
R6575 VSS.n2600 VSS.n254 40.8246
R6576 VSS.n2595 VSS.n253 40.8246
R6577 VSS.n1500 VSS.n286 40.8246
R6578 VSS.n1505 VSS.n287 40.8246
R6579 VSS.n1510 VSS.n288 40.8246
R6580 VSS.n1515 VSS.n289 40.8246
R6581 VSS.n1561 VSS.n1559 40.8246
R6582 VSS.n1658 VSS.n1657 40.8246
R6583 VSS.n1660 VSS.n1659 40.8246
R6584 VSS.n1663 VSS.n1656 40.8246
R6585 VSS.n1665 VSS.n1664 40.8246
R6586 VSS.n1667 VSS.n1666 40.8246
R6587 VSS.n1670 VSS.n1654 40.8246
R6588 VSS.n1672 VSS.n1671 40.8246
R6589 VSS.n1674 VSS.n1673 40.8246
R6590 VSS.n1677 VSS.n1652 40.8246
R6591 VSS.n1678 VSS.n1677 40.8246
R6592 VSS.n1651 VSS.n1614 40.8246
R6593 VSS.n1649 VSS.n1648 40.8246
R6594 VSS.n1647 VSS.n1646 40.8246
R6595 VSS.n1645 VSS.n1644 40.8246
R6596 VSS.n1641 VSS.n1616 40.8246
R6597 VSS.n1640 VSS.n1639 40.8246
R6598 VSS.n1638 VSS.n1637 40.8246
R6599 VSS.n1636 VSS.n1635 40.8246
R6600 VSS.n1632 VSS.n1619 40.8246
R6601 VSS.n1631 VSS.n1630 40.8246
R6602 VSS.n1629 VSS.n1628 40.8246
R6603 VSS.n1627 VSS.n1626 40.8246
R6604 VSS.n1623 VSS.n1622 40.8246
R6605 VSS.n5220 VSS.n5219 40.8246
R6606 VSS.n5218 VSS.n5217 40.8246
R6607 VSS.n5216 VSS.n5215 40.8246
R6608 VSS.n5212 VSS.n409 40.8246
R6609 VSS.n5211 VSS.n5210 40.8246
R6610 VSS.n5209 VSS.n5208 40.8246
R6611 VSS.n5207 VSS.n5206 40.8246
R6612 VSS.n5203 VSS.n412 40.8246
R6613 VSS.n5202 VSS.n5201 40.8246
R6614 VSS.n5200 VSS.n5199 40.8246
R6615 VSS.n5199 VSS.n414 40.8246
R6616 VSS.n5194 VSS.n417 40.8246
R6617 VSS.n5192 VSS.n418 40.8246
R6618 VSS.n1363 VSS.n1362 40.8246
R6619 VSS.n1366 VSS.n1364 40.8246
R6620 VSS.n1368 VSS.n1367 40.8246
R6621 VSS.n1370 VSS.n1369 40.8246
R6622 VSS.n1373 VSS.n1360 40.8246
R6623 VSS.n1375 VSS.n1374 40.8246
R6624 VSS.n1377 VSS.n1376 40.8246
R6625 VSS.n1380 VSS.n1358 40.8246
R6626 VSS.n1382 VSS.n1381 40.8246
R6627 VSS.n1383 VSS.n1382 40.8246
R6628 VSS.n1387 VSS.n1356 40.8246
R6629 VSS.n3214 VSS.n3213 40.8246
R6630 VSS.n3212 VSS.n3211 40.8246
R6631 VSS.n3210 VSS.n3209 40.8246
R6632 VSS.n3206 VSS.n3181 40.8246
R6633 VSS.n3205 VSS.n3204 40.8246
R6634 VSS.n3203 VSS.n3202 40.8246
R6635 VSS.n3201 VSS.n3200 40.8246
R6636 VSS.n3197 VSS.n3184 40.8246
R6637 VSS.n3196 VSS.n3195 40.8246
R6638 VSS.n3194 VSS.n3193 40.8246
R6639 VSS.n3192 VSS.n3191 40.8246
R6640 VSS.n3188 VSS.n3187 40.8246
R6641 VSS.n4473 VSS.n4471 40.8246
R6642 VSS.n4475 VSS.n4474 40.8246
R6643 VSS.n4477 VSS.n4476 40.8246
R6644 VSS.n4480 VSS.n4468 40.8246
R6645 VSS.n4482 VSS.n4481 40.8246
R6646 VSS.n4484 VSS.n4483 40.8246
R6647 VSS.n4487 VSS.n4466 40.8246
R6648 VSS.n4489 VSS.n4488 40.8246
R6649 VSS.n4491 VSS.n4490 40.8246
R6650 VSS.n4495 VSS.n4464 40.8246
R6651 VSS.n4496 VSS.n4495 40.8246
R6652 VSS.n4499 VSS.n4498 40.8246
R6653 VSS.n4491 VSS.n4464 40.8246
R6654 VSS.n4488 VSS.n4487 40.8246
R6655 VSS.n4483 VSS.n4482 40.8246
R6656 VSS.n4477 VSS.n4468 40.8246
R6657 VSS.n4474 VSS.n4473 40.8246
R6658 VSS.n3191 VSS.n3187 40.8246
R6659 VSS.n3195 VSS.n3194 40.8246
R6660 VSS.n3200 VSS.n3184 40.8246
R6661 VSS.n3204 VSS.n3203 40.8246
R6662 VSS.n3209 VSS.n3181 40.8246
R6663 VSS.n3213 VSS.n3212 40.8246
R6664 VSS.n5201 VSS.n5200 40.8246
R6665 VSS.n5206 VSS.n412 40.8246
R6666 VSS.n5210 VSS.n5209 40.8246
R6667 VSS.n5215 VSS.n409 40.8246
R6668 VSS.n5219 VSS.n5218 40.8246
R6669 VSS.n1626 VSS.n1622 40.8246
R6670 VSS.n1630 VSS.n1629 40.8246
R6671 VSS.n1635 VSS.n1619 40.8246
R6672 VSS.n1639 VSS.n1638 40.8246
R6673 VSS.n1644 VSS.n1616 40.8246
R6674 VSS.n1674 VSS.n1652 40.8246
R6675 VSS.n1671 VSS.n1670 40.8246
R6676 VSS.n1666 VSS.n1665 40.8246
R6677 VSS.n1660 VSS.n1656 40.8246
R6678 VSS.n1657 VSS.n1561 40.8246
R6679 VSS.n2530 VSS.n1559 40.8246
R6680 VSS.n4490 VSS.n4489 40.8246
R6681 VSS.n4484 VSS.n4466 40.8246
R6682 VSS.n4481 VSS.n4480 40.8246
R6683 VSS.n4476 VSS.n4475 40.8246
R6684 VSS.n4471 VSS.n4470 40.8246
R6685 VSS.n3193 VSS.n3192 40.8246
R6686 VSS.n3197 VSS.n3196 40.8246
R6687 VSS.n3202 VSS.n3201 40.8246
R6688 VSS.n3206 VSS.n3205 40.8246
R6689 VSS.n3211 VSS.n3210 40.8246
R6690 VSS.n5203 VSS.n5202 40.8246
R6691 VSS.n5208 VSS.n5207 40.8246
R6692 VSS.n5212 VSS.n5211 40.8246
R6693 VSS.n5217 VSS.n5216 40.8246
R6694 VSS.n5221 VSS.n5220 40.8246
R6695 VSS.n1628 VSS.n1627 40.8246
R6696 VSS.n1632 VSS.n1631 40.8246
R6697 VSS.n1637 VSS.n1636 40.8246
R6698 VSS.n1641 VSS.n1640 40.8246
R6699 VSS.n1646 VSS.n1645 40.8246
R6700 VSS.n1673 VSS.n1672 40.8246
R6701 VSS.n1667 VSS.n1654 40.8246
R6702 VSS.n1664 VSS.n1663 40.8246
R6703 VSS.n1659 VSS.n1658 40.8246
R6704 VSS.n1377 VSS.n1358 40.8246
R6705 VSS.n1374 VSS.n1373 40.8246
R6706 VSS.n1369 VSS.n1368 40.8246
R6707 VSS.n1364 VSS.n1363 40.8246
R6708 VSS.n1381 VSS.n1380 40.8246
R6709 VSS.n1376 VSS.n1375 40.8246
R6710 VSS.n1370 VSS.n1360 40.8246
R6711 VSS.n1367 VSS.n1366 40.8246
R6712 VSS.n1384 VSS.n1383 40.8246
R6713 VSS.n3215 VSS.n3214 40.8246
R6714 VSS.n1384 VSS.n1356 40.8246
R6715 VSS.n3220 VSS.n3219 40.8246
R6716 VSS.n497 VSS.n496 40.8246
R6717 VSS.n492 VSS.n491 40.8246
R6718 VSS.n490 VSS.n489 40.8246
R6719 VSS.n488 VSS.n487 40.8246
R6720 VSS.n5147 VSS.n457 40.8246
R6721 VSS.n5149 VSS.n5148 40.8246
R6722 VSS.n5151 VSS.n5150 40.8246
R6723 VSS.n3217 VSS.n453 40.8246
R6724 VSS.n4879 VSS.n4878 40.8246
R6725 VSS.n4871 VSS.n504 40.8246
R6726 VSS.n4870 VSS.n4869 40.8246
R6727 VSS.n4862 VSS.n505 40.8246
R6728 VSS.n4861 VSS.n4860 40.8246
R6729 VSS.n4849 VSS.n506 40.8246
R6730 VSS.n4848 VSS.n4847 40.8246
R6731 VSS.n514 VSS.n507 40.8246
R6732 VSS.n5118 VSS.n509 40.8246
R6733 VSS.n5119 VSS.n508 40.8246
R6734 VSS.n5124 VSS.n5123 40.8246
R6735 VSS.n681 VSS.n680 40.8246
R6736 VSS.n1893 VSS.n1889 40.8246
R6737 VSS.n1894 VSS.n1893 40.8246
R6738 VSS.n5121 VSS.n502 40.8246
R6739 VSS.n703 VSS.n684 40.8246
R6740 VSS.n700 VSS.n699 40.8246
R6741 VSS.n695 VSS.n694 40.8246
R6742 VSS.n690 VSS.n689 40.8246
R6743 VSS.n701 VSS.n679 40.8246
R6744 VSS.n696 VSS.n678 40.8246
R6745 VSS.n691 VSS.n677 40.8246
R6746 VSS.n686 VSS.n676 40.8246
R6747 VSS.n4557 VSS.n671 40.8246
R6748 VSS.n4680 VSS.n711 40.8246
R6749 VSS.n683 VSS.n682 40.8246
R6750 VSS.n4682 VSS.n4681 40.8246
R6751 VSS.n709 VSS.n683 40.8246
R6752 VSS.n4780 VSS.n4684 40.8246
R6753 VSS.n4777 VSS.n4691 40.8246
R6754 VSS.n4778 VSS.n4690 40.8246
R6755 VSS.n4733 VSS.n4732 40.8246
R6756 VSS.n4735 VSS.n4689 40.8246
R6757 VSS.n4736 VSS.n4734 40.8246
R6758 VSS.n4738 VSS.n4688 40.8246
R6759 VSS.n4739 VSS.n4737 40.8246
R6760 VSS.n4742 VSS.n4687 40.8246
R6761 VSS.n4741 VSS.n4731 40.8246
R6762 VSS.n4686 VSS.n4685 40.8246
R6763 VSS.n3896 VSS.n3895 40.8246
R6764 VSS.n3895 VSS.n272 40.8246
R6765 VSS.n4498 VSS.n4497 40.8246
R6766 VSS.n4497 VSS.n4496 40.8246
R6767 VSS.n4657 VSS.n719 40.8246
R6768 VSS.n4658 VSS.n4657 40.8246
R6769 VSS.n3758 VSS.n3757 40.8246
R6770 VSS.n3759 VSS.n3581 40.8246
R6771 VSS.n3656 VSS.n3655 40.8246
R6772 VSS.n3656 VSS.n3585 40.8246
R6773 VSS.n3665 VSS.n3664 40.8246
R6774 VSS.n3665 VSS.n3586 40.8246
R6775 VSS.n3674 VSS.n3673 40.8246
R6776 VSS.n3674 VSS.n3587 40.8246
R6777 VSS.n3708 VSS.n3707 40.8246
R6778 VSS.n3584 VSS.n960 40.8246
R6779 VSS.n1009 VSS.n964 40.8246
R6780 VSS.n1010 VSS.n964 40.8246
R6781 VSS.n4206 VSS.n965 40.8246
R6782 VSS.n4207 VSS.n4206 40.8246
R6783 VSS.n4211 VSS.n966 40.8246
R6784 VSS.n4212 VSS.n4211 40.8246
R6785 VSS.n4216 VSS.n967 40.8246
R6786 VSS.n4217 VSS.n4216 40.8246
R6787 VSS.n4221 VSS.n968 40.8246
R6788 VSS.n4222 VSS.n4221 40.8246
R6789 VSS.n4201 VSS.n969 40.8246
R6790 VSS.n4202 VSS.n1005 40.8246
R6791 VSS.n4204 VSS.n4203 40.8246
R6792 VSS.n4250 VSS.n971 40.8246
R6793 VSS.n4250 VSS.n4249 40.8246
R6794 VSS.n4245 VSS.n972 40.8246
R6795 VSS.n4245 VSS.n4244 40.8246
R6796 VSS.n4240 VSS.n973 40.8246
R6797 VSS.n4240 VSS.n4239 40.8246
R6798 VSS.n4235 VSS.n974 40.8246
R6799 VSS.n4235 VSS.n4234 40.8246
R6800 VSS.n4230 VSS.n975 40.8246
R6801 VSS.n4230 VSS.n4229 40.8246
R6802 VSS.n4225 VSS.n976 40.8246
R6803 VSS.n3309 VSS.n977 40.8246
R6804 VSS.n3310 VSS.n3309 40.8246
R6805 VSS.n3314 VSS.n978 40.8246
R6806 VSS.n3315 VSS.n3314 40.8246
R6807 VSS.n3319 VSS.n979 40.8246
R6808 VSS.n3320 VSS.n3319 40.8246
R6809 VSS.n3324 VSS.n980 40.8246
R6810 VSS.n3325 VSS.n3324 40.8246
R6811 VSS.n3329 VSS.n981 40.8246
R6812 VSS.n3330 VSS.n3329 40.8246
R6813 VSS.n3339 VSS.n982 40.8246
R6814 VSS.n3338 VSS.n1004 40.8246
R6815 VSS.n3336 VSS.n3334 40.8246
R6816 VSS.n3306 VSS.n984 40.8246
R6817 VSS.n3306 VSS.n3305 40.8246
R6818 VSS.n3301 VSS.n985 40.8246
R6819 VSS.n3301 VSS.n3300 40.8246
R6820 VSS.n3296 VSS.n986 40.8246
R6821 VSS.n3296 VSS.n3295 40.8246
R6822 VSS.n3291 VSS.n987 40.8246
R6823 VSS.n3291 VSS.n3290 40.8246
R6824 VSS.n3286 VSS.n988 40.8246
R6825 VSS.n3286 VSS.n3285 40.8246
R6826 VSS.n3281 VSS.n989 40.8246
R6827 VSS.n3829 VSS.n990 40.8246
R6828 VSS.n3829 VSS.n3828 40.8246
R6829 VSS.n3824 VSS.n991 40.8246
R6830 VSS.n3824 VSS.n3823 40.8246
R6831 VSS.n3819 VSS.n992 40.8246
R6832 VSS.n3819 VSS.n3818 40.8246
R6833 VSS.n3814 VSS.n993 40.8246
R6834 VSS.n3814 VSS.n3813 40.8246
R6835 VSS.n3809 VSS.n994 40.8246
R6836 VSS.n3809 VSS.n3808 40.8246
R6837 VSS.n3804 VSS.n995 40.8246
R6838 VSS.n3804 VSS.n3803 40.8246
R6839 VSS.n4401 VSS.n962 40.8246
R6840 VSS.n1246 VSS.n997 40.8246
R6841 VSS.n1247 VSS.n1246 40.8246
R6842 VSS.n1251 VSS.n998 40.8246
R6843 VSS.n1252 VSS.n1251 40.8246
R6844 VSS.n1256 VSS.n999 40.8246
R6845 VSS.n1257 VSS.n1256 40.8246
R6846 VSS.n1261 VSS.n1000 40.8246
R6847 VSS.n1262 VSS.n1261 40.8246
R6848 VSS.n1266 VSS.n1001 40.8246
R6849 VSS.n1266 VSS.n1265 40.8246
R6850 VSS.n3960 VSS.n1243 40.8246
R6851 VSS.n4022 VSS.n1117 40.8246
R6852 VSS.n4022 VSS.n4021 40.8246
R6853 VSS.n3795 VSS.n3794 40.8246
R6854 VSS.n3794 VSS.n1119 40.8246
R6855 VSS.n3531 VSS.n3526 40.8246
R6856 VSS.n3531 VSS.n1120 40.8246
R6857 VSS.n3572 VSS.n3525 40.8246
R6858 VSS.n3572 VSS.n1121 40.8246
R6859 VSS.n3564 VSS.n3524 40.8246
R6860 VSS.n3564 VSS.n1122 40.8246
R6861 VSS.n3797 VSS.n1123 40.8246
R6862 VSS.n4019 VSS.n1117 40.8246
R6863 VSS.n3707 VSS.n3584 40.8246
R6864 VSS.n3709 VSS.n3708 40.8246
R6865 VSS.n3588 VSS.n3587 40.8246
R6866 VSS.n3672 VSS.n3586 40.8246
R6867 VSS.n3673 VSS.n3672 40.8246
R6868 VSS.n3663 VSS.n3585 40.8246
R6869 VSS.n3664 VSS.n3663 40.8246
R6870 VSS.n3654 VSS.n3581 40.8246
R6871 VSS.n3655 VSS.n3654 40.8246
R6872 VSS.n3759 VSS.n3758 40.8246
R6873 VSS.n3798 VSS.n1122 40.8246
R6874 VSS.n3798 VSS.n3797 40.8246
R6875 VSS.n3560 VSS.n1121 40.8246
R6876 VSS.n3560 VSS.n3524 40.8246
R6877 VSS.n3552 VSS.n1120 40.8246
R6878 VSS.n3552 VSS.n3525 40.8246
R6879 VSS.n3529 VSS.n1119 40.8246
R6880 VSS.n3529 VSS.n3526 40.8246
R6881 VSS.n4021 VSS.n1118 40.8246
R6882 VSS.n3795 VSS.n1118 40.8246
R6883 VSS.n5456 VSS.n77 40.8246
R6884 VSS.n5454 VSS.n5453 40.8246
R6885 VSS.n5453 VSS.n78 40.8246
R6886 VSS.n120 VSS.n116 40.8246
R6887 VSS.n120 VSS.n79 40.8246
R6888 VSS.n125 VSS.n115 40.8246
R6889 VSS.n125 VSS.n80 40.8246
R6890 VSS.n88 VSS.n83 40.8246
R6891 VSS.n88 VSS.n81 40.8246
R6892 VSS.n82 VSS.n75 40.8246
R6893 VSS.n5472 VSS.n82 40.8246
R6894 VSS.n2894 VSS.n250 40.8246
R6895 VSS.n5373 VSS.n245 40.8246
R6896 VSS.n259 VSS.n258 40.8246
R6897 VSS.n260 VSS.n259 40.8246
R6898 VSS.n5193 VSS.n5192 40.8246
R6899 VSS.n5195 VSS.n5194 40.8246
R6900 VSS.n1362 VSS.n418 40.8246
R6901 VSS.n5195 VSS.n414 40.8246
R6902 VSS.n1876 VSS.n1875 40.8246
R6903 VSS.n1872 VSS.n423 40.8246
R6904 VSS.n1873 VSS.n1814 40.8246
R6905 VSS.n1837 VSS.n424 40.8246
R6906 VSS.n1828 VSS.n1813 40.8246
R6907 VSS.n1824 VSS.n425 40.8246
R6908 VSS.n1812 VSS.n1811 40.8246
R6909 VSS.n433 VSS.n426 40.8246
R6910 VSS.n5187 VSS.n428 40.8246
R6911 VSS.n5188 VSS.n427 40.8246
R6912 VSS.n5190 VSS.n421 40.8246
R6913 VSS.n1915 VSS.n1914 40.8246
R6914 VSS.n1919 VSS.n1879 40.8246
R6915 VSS.n1951 VSS.n1878 40.8246
R6916 VSS.n1951 VSS.n1950 40.8246
R6917 VSS.n4949 VSS.n629 40.8246
R6918 VSS.n4946 VSS.n4945 40.8246
R6919 VSS.n4947 VSS.n634 40.8246
R6920 VSS.n4910 VSS.n4909 40.8246
R6921 VSS.n4918 VSS.n633 40.8246
R6922 VSS.n4917 VSS.n4916 40.8246
R6923 VSS.n4929 VSS.n632 40.8246
R6924 VSS.n4931 VSS.n4930 40.8246
R6925 VSS.n661 VSS.n631 40.8246
R6926 VSS.n660 VSS.n659 40.8246
R6927 VSS.n1917 VSS.n630 40.8246
R6928 VSS.n1107 VSS.n1106 40.8246
R6929 VSS.n1106 VSS.n1105 40.8246
R6930 VSS.n1072 VSS.n1066 40.8246
R6931 VSS.n1072 VSS.n1067 40.8246
R6932 VSS.n1089 VSS.n1065 40.8246
R6933 VSS.n1090 VSS.n1089 40.8246
R6934 VSS.n4146 VSS.n1064 40.8246
R6935 VSS.n1081 VSS.n1064 40.8246
R6936 VSS.n4149 VSS.n1062 40.8246
R6937 VSS.n4149 VSS.n4148 40.8246
R6938 VSS.n4143 VSS.n4142 40.8246
R6939 VSS.n4308 VSS.n4255 40.8246
R6940 VSS.n4306 VSS.n4305 40.8246
R6941 VSS.n4305 VSS.n4200 40.8246
R6942 VSS.n4268 VSS.n4259 40.8246
R6943 VSS.n4269 VSS.n4268 40.8246
R6944 VSS.n4270 VSS.n4258 40.8246
R6945 VSS.n4272 VSS.n4270 40.8246
R6946 VSS.n4279 VSS.n4257 40.8246
R6947 VSS.n4279 VSS.n4278 40.8246
R6948 VSS.n4273 VSS.n4256 40.8246
R6949 VSS.n4275 VSS.n4273 40.8246
R6950 VSS.n2594 VSS.n249 40.8246
R6951 VSS.n5371 VSS.n292 40.8246
R6952 VSS.n5369 VSS.n5368 40.8246
R6953 VSS.n5369 VSS.n252 40.8246
R6954 VSS.n1648 VSS.n1647 40.8246
R6955 VSS.n1650 VSS.n1649 40.8246
R6956 VSS.n1679 VSS.n1651 40.8246
R6957 VSS.n1679 VSS.n1678 40.8246
R6958 VSS.n2472 VSS.n1698 40.8246
R6959 VSS.n2474 VSS.n2473 40.8246
R6960 VSS.n2476 VSS.n2475 40.8246
R6961 VSS.n1693 VSS.n1612 40.8246
R6962 VSS.n1694 VSS.n1689 40.8246
R6963 VSS.n1688 VSS.n1687 40.8246
R6964 VSS.n2492 VSS.n1585 40.8246
R6965 VSS.n2494 VSS.n2493 40.8246
R6966 VSS.n1683 VSS.n1583 40.8246
R6967 VSS.n1685 VSS.n1684 40.8246
R6968 VSS.n1686 VSS.n1682 40.8246
R6969 VSS.n2167 VSS.n2166 40.8246
R6970 VSS.n2165 VSS.n1999 40.8246
R6971 VSS.n2162 VSS.n2161 40.8246
R6972 VSS.n2163 VSS.n2162 40.8246
R6973 VSS.n2359 VSS.n2358 40.8246
R6974 VSS.n2355 VSS.n2069 40.8246
R6975 VSS.n2356 VSS.n2075 40.8246
R6976 VSS.n2099 VSS.n2098 40.8246
R6977 VSS.n2090 VSS.n2074 40.8246
R6978 VSS.n2089 VSS.n2088 40.8246
R6979 VSS.n2073 VSS.n2072 40.8246
R6980 VSS.n2071 VSS.n2070 40.8246
R6981 VSS.n2460 VSS.n2005 40.8246
R6982 VSS.n2462 VSS.n2461 40.8246
R6983 VSS.n2466 VSS.n2000 40.8246
R6984 VSS.n324 VSS.n296 40.8246
R6985 VSS.n5317 VSS.n297 40.8246
R6986 VSS.n5318 VSS.n322 40.8246
R6987 VSS.n2692 VSS.n298 40.8246
R6988 VSS.n2682 VSS.n321 40.8246
R6989 VSS.n5321 VSS.n299 40.8246
R6990 VSS.n5320 VSS.n316 40.8246
R6991 VSS.n319 VSS.n300 40.8246
R6992 VSS.n320 VSS.n318 40.8246
R6993 VSS.n5359 VSS.n301 40.8246
R6994 VSS.n5363 VSS.n303 40.8246
R6995 VSS.n2725 VSS.n2724 40.8246
R6996 VSS.n2721 VSS.n155 40.8246
R6997 VSS.n2722 VSS.n2643 40.8246
R6998 VSS.n2663 VSS.n156 40.8246
R6999 VSS.n2654 VSS.n2642 40.8246
R7000 VSS.n2652 VSS.n157 40.8246
R7001 VSS.n2641 VSS.n2640 40.8246
R7002 VSS.n167 VSS.n158 40.8246
R7003 VSS.n5423 VSS.n160 40.8246
R7004 VSS.n5424 VSS.n159 40.8246
R7005 VSS.n5426 VSS.n153 40.8246
R7006 VSS.n5379 VSS.n234 40.8246
R7007 VSS.n5381 VSS.n5380 40.8246
R7008 VSS.n5389 VSS.n231 40.8246
R7009 VSS.n5391 VSS.n5390 40.8246
R7010 VSS.n230 VSS.n229 40.8246
R7011 VSS.n222 VSS.n221 40.8246
R7012 VSS.n5403 VSS.n199 40.8246
R7013 VSS.n5405 VSS.n5404 40.8246
R7014 VSS.n3343 VSS.n197 40.8246
R7015 VSS.n3345 VSS.n3344 40.8246
R7016 VSS.n3347 VSS.n3346 40.8246
R7017 VSS.n3838 VSS.n3837 40.8246
R7018 VSS.n3392 VSS.n1343 40.8246
R7019 VSS.n3394 VSS.n3393 40.8246
R7020 VSS.n3383 VSS.n3257 40.8246
R7021 VSS.n3382 VSS.n3381 40.8246
R7022 VSS.n3408 VSS.n3258 40.8246
R7023 VSS.n3410 VSS.n3409 40.8246
R7024 VSS.n3371 VSS.n3259 40.8246
R7025 VSS.n3370 VSS.n3369 40.8246
R7026 VSS.n3504 VSS.n3260 40.8246
R7027 VSS.n3834 VSS.n3262 40.8246
R7028 VSS.n1304 VSS.n948 40.8246
R7029 VSS.n3870 VSS.n951 40.8246
R7030 VSS.n3869 VSS.n1310 40.8246
R7031 VSS.n3866 VSS.n952 40.8246
R7032 VSS.n3867 VSS.n1313 40.8246
R7033 VSS.n3454 VSS.n953 40.8246
R7034 VSS.n3450 VSS.n1312 40.8246
R7035 VSS.n3472 VSS.n954 40.8246
R7036 VSS.n3422 VSS.n1311 40.8246
R7037 VSS.n3420 VSS.n955 40.8246
R7038 VSS.n4404 VSS.n957 40.8246
R7039 VSS.n1243 VSS.n1002 40.8246
R7040 VSS.n1265 VSS.n1002 40.8246
R7041 VSS.n1263 VSS.n1262 40.8246
R7042 VSS.n1258 VSS.n1257 40.8246
R7043 VSS.n1253 VSS.n1252 40.8246
R7044 VSS.n1248 VSS.n1247 40.8246
R7045 VSS.n996 VSS.n962 40.8246
R7046 VSS.n3803 VSS.n1003 40.8246
R7047 VSS.n3808 VSS.n3807 40.8246
R7048 VSS.n3813 VSS.n3812 40.8246
R7049 VSS.n3818 VSS.n3817 40.8246
R7050 VSS.n3823 VSS.n3822 40.8246
R7051 VSS.n3828 VSS.n3827 40.8246
R7052 VSS.n3285 VSS.n3284 40.8246
R7053 VSS.n3290 VSS.n3289 40.8246
R7054 VSS.n3295 VSS.n3294 40.8246
R7055 VSS.n3300 VSS.n3299 40.8246
R7056 VSS.n3305 VSS.n3304 40.8246
R7057 VSS.n3336 VSS.n983 40.8246
R7058 VSS.n3339 VSS.n3338 40.8246
R7059 VSS.n3331 VSS.n3330 40.8246
R7060 VSS.n3326 VSS.n3325 40.8246
R7061 VSS.n3321 VSS.n3320 40.8246
R7062 VSS.n3316 VSS.n3315 40.8246
R7063 VSS.n3311 VSS.n3310 40.8246
R7064 VSS.n4229 VSS.n4228 40.8246
R7065 VSS.n4234 VSS.n4233 40.8246
R7066 VSS.n4239 VSS.n4238 40.8246
R7067 VSS.n4244 VSS.n4243 40.8246
R7068 VSS.n4249 VSS.n4248 40.8246
R7069 VSS.n4204 VSS.n970 40.8246
R7070 VSS.n4202 VSS.n4201 40.8246
R7071 VSS.n4223 VSS.n4222 40.8246
R7072 VSS.n4218 VSS.n4217 40.8246
R7073 VSS.n4213 VSS.n4212 40.8246
R7074 VSS.n4208 VSS.n4207 40.8246
R7075 VSS.n1011 VSS.n1010 40.8246
R7076 VSS.n4399 VSS.n1009 40.8246
R7077 VSS.n1263 VSS.n1001 40.8246
R7078 VSS.n1258 VSS.n1000 40.8246
R7079 VSS.n1253 VSS.n999 40.8246
R7080 VSS.n1248 VSS.n998 40.8246
R7081 VSS.n997 VSS.n996 40.8246
R7082 VSS.n3807 VSS.n995 40.8246
R7083 VSS.n3812 VSS.n994 40.8246
R7084 VSS.n3817 VSS.n993 40.8246
R7085 VSS.n3822 VSS.n992 40.8246
R7086 VSS.n3827 VSS.n991 40.8246
R7087 VSS.n3831 VSS.n990 40.8246
R7088 VSS.n3284 VSS.n989 40.8246
R7089 VSS.n3289 VSS.n988 40.8246
R7090 VSS.n3294 VSS.n987 40.8246
R7091 VSS.n3299 VSS.n986 40.8246
R7092 VSS.n3304 VSS.n985 40.8246
R7093 VSS.n3334 VSS.n984 40.8246
R7094 VSS.n3331 VSS.n982 40.8246
R7095 VSS.n3326 VSS.n981 40.8246
R7096 VSS.n3321 VSS.n980 40.8246
R7097 VSS.n3316 VSS.n979 40.8246
R7098 VSS.n3311 VSS.n978 40.8246
R7099 VSS.n1007 VSS.n977 40.8246
R7100 VSS.n4228 VSS.n976 40.8246
R7101 VSS.n4233 VSS.n975 40.8246
R7102 VSS.n4238 VSS.n974 40.8246
R7103 VSS.n4243 VSS.n973 40.8246
R7104 VSS.n4248 VSS.n972 40.8246
R7105 VSS.n4203 VSS.n971 40.8246
R7106 VSS.n4223 VSS.n969 40.8246
R7107 VSS.n4218 VSS.n968 40.8246
R7108 VSS.n4213 VSS.n967 40.8246
R7109 VSS.n4208 VSS.n966 40.8246
R7110 VSS.n1011 VSS.n965 40.8246
R7111 VSS.t31 VSS.n1129 40.6176
R7112 VSS.n5558 VSS.t14 40.0612
R7113 VSS.t16 VSS.n1138 40.0612
R7114 VSS.n5528 VSS.t93 39.5048
R7115 VSS.n68 VSS.t25 38.392
R7116 VSS.t3 VSS.n69 38.392
R7117 VSS.n4013 VSS.n4012 36.563
R7118 VSS.n4014 VSS.n4013 36.563
R7119 VSS.n1163 VSS.n1162 36.563
R7120 VSS.n1162 VSS.n1161 36.563
R7121 VSS.n58 VSS.n57 36.563
R7122 VSS.n3722 VSS.n58 36.563
R7123 VSS.n5504 VSS.n5503 36.563
R7124 VSS.n5503 VSS.n5502 36.563
R7125 VSS.t10 VSS.n5563 35.61
R7126 VSS.t32 VSS.t42 35.0536
R7127 VSS.n1173 VSS.n1169 34.4123
R7128 VSS.n1169 VSS.n1168 34.4123
R7129 VSS.n1182 VSS.n1181 34.4123
R7130 VSS.n1183 VSS.n1182 34.4123
R7131 VSS.t54 VSS.n14 33.9408
R7132 VSS.n5527 VSS.t54 33.9408
R7133 VSS.t54 VSS.n68 33.9408
R7134 VSS.n1160 VSS.t54 33.9408
R7135 VSS.t54 VSS.n3734 33.9408
R7136 VSS.n5508 VSS.n49 33.9393
R7137 VSS.t39 VSS.n1152 33.3844
R7138 VSS.n3725 VSS.n3722 32.2716
R7139 VSS.n26 VSS.n25 30.79
R7140 VSS.t26 VSS.n5494 30.6024
R7141 VSS.n5478 VSS.t5 30.6024
R7142 VSS.n674 VSS.n345 30.0246
R7143 VSS.n247 VSS.n244 30.0246
R7144 VSS.n406 VSS.n343 30.0246
R7145 VSS.n1008 VSS.n963 30.0246
R7146 VSS.n710 VSS.n345 29.4359
R7147 VSS.n5372 VSS.n247 29.4359
R7148 VSS.n407 VSS.n343 29.4359
R7149 VSS.n4400 VSS.n963 29.4359
R7150 VSS.n1154 VSS.t4 28.9332
R7151 VSS.n1147 VSS.t45 28.9332
R7152 VSS.n5556 VSS.t65 27.8204
R7153 VSS.n1161 VSS.t105 27.8204
R7154 VSS.n5501 VSS.t19 27.264
R7155 VSS.n1154 VSS.t6 25.5948
R7156 VSS.t6 VSS.n1145 24.482
R7157 VSS.n4651 VSS.n720 24.3817
R7158 VSS.n3894 VSS.n897 24.3817
R7159 VSS.n4499 VSS.n784 24.3817
R7160 VSS.n3960 VSS.n1244 24.3817
R7161 VSS.n1180 VSS.t9 23.1325
R7162 VSS.n1170 VSS.t8 23.0375
R7163 VSS.n64 VSS.t19 22.8128
R7164 VSS.n14 VSS.t65 22.2564
R7165 VSS.n1178 VSS.t38 21.5736
R7166 VSS.n1171 VSS.t2 21.5494
R7167 VSS.n1171 VSS.t37 21.4809
R7168 VSS.t4 VSS.n1153 21.1436
R7169 VSS.n1152 VSS.t45 21.1436
R7170 VSS.n5509 VSS.n0 20.5168
R7171 VSS.n5567 VSS.n5566 20.0506
R7172 VSS.n5511 VSS.t17 20.0308
R7173 VSS.n1191 VSS.n49 19.8035
R7174 VSS.n5495 VSS.t26 19.4745
R7175 VSS.t5 VSS.n5477 19.4745
R7176 VSS.n5502 VSS.n59 18.9181
R7177 VSS.t105 VSS.n1160 17.8053
R7178 VSS.n5512 VSS.n5511 17.2489
R7179 VSS.n5044 VSS.n594 17.1965
R7180 VSS.n1153 VSS.t39 16.6925
R7181 VSS.n3997 VSS.n1199 16.6357
R7182 VSS.n5550 VSS.t54 16.1361
R7183 VSS.t54 VSS.n5526 16.1361
R7184 VSS.n5487 VSS.t54 16.1361
R7185 VSS.n3736 VSS.t54 16.1361
R7186 VSS.n4180 VSS.n4179 16.0005
R7187 VSS.n4179 VSS.n4178 16.0005
R7188 VSS.n4178 VSS.n4176 16.0005
R7189 VSS.n4176 VSS.n4173 16.0005
R7190 VSS.n4173 VSS.n4172 16.0005
R7191 VSS.n4172 VSS.n4169 16.0005
R7192 VSS.n4169 VSS.n4168 16.0005
R7193 VSS.n4168 VSS.n146 16.0005
R7194 VSS.n5431 VSS.n5430 16.0005
R7195 VSS.n5431 VSS.n144 16.0005
R7196 VSS.n5437 VSS.n144 16.0005
R7197 VSS.n5438 VSS.n5437 16.0005
R7198 VSS.n5439 VSS.n5438 16.0005
R7199 VSS.n5439 VSS.n142 16.0005
R7200 VSS.n5444 VSS.n142 16.0005
R7201 VSS.n5445 VSS.n5444 16.0005
R7202 VSS.n3508 VSS.n3507 16.0005
R7203 VSS.n3510 VSS.n3508 16.0005
R7204 VSS.n3511 VSS.n3510 16.0005
R7205 VSS.n3514 VSS.n3511 16.0005
R7206 VSS.n3515 VSS.n3514 16.0005
R7207 VSS.n3518 VSS.n3515 16.0005
R7208 VSS.n3520 VSS.n3518 16.0005
R7209 VSS.n3521 VSS.n3520 16.0005
R7210 VSS.n3592 VSS.n3522 16.0005
R7211 VSS.n3593 VSS.n3592 16.0005
R7212 VSS.n3596 VSS.n3593 16.0005
R7213 VSS.n3597 VSS.n3596 16.0005
R7214 VSS.n3600 VSS.n3597 16.0005
R7215 VSS.n3601 VSS.n3600 16.0005
R7216 VSS.n3604 VSS.n3601 16.0005
R7217 VSS.n3608 VSS.n3604 16.0005
R7218 VSS.n3775 VSS.n1114 16.0005
R7219 VSS.n3775 VSS.n3774 16.0005
R7220 VSS.n3774 VSS.n3771 16.0005
R7221 VSS.n3771 VSS.n3770 16.0005
R7222 VSS.n3770 VSS.n3768 16.0005
R7223 VSS.n3768 VSS.n3767 16.0005
R7224 VSS.n3767 VSS.n3765 16.0005
R7225 VSS.n3765 VSS.n3762 16.0005
R7226 VSS.n3636 VSS.n3578 16.0005
R7227 VSS.n3636 VSS.n3635 16.0005
R7228 VSS.n3635 VSS.n3634 16.0005
R7229 VSS.n3634 VSS.n3618 16.0005
R7230 VSS.n3629 VSS.n3618 16.0005
R7231 VSS.n3629 VSS.n3628 16.0005
R7232 VSS.n3628 VSS.n3627 16.0005
R7233 VSS.n3627 VSS.n1216 16.0005
R7234 VSS.n3704 VSS.n3609 16.0005
R7235 VSS.n3699 VSS.n3609 16.0005
R7236 VSS.n3699 VSS.n3698 16.0005
R7237 VSS.n3698 VSS.n3697 16.0005
R7238 VSS.n3697 VSS.n3686 16.0005
R7239 VSS.n3692 VSS.n3686 16.0005
R7240 VSS.n3692 VSS.n3691 16.0005
R7241 VSS.n3691 VSS.n3690 16.0005
R7242 VSS.n3443 VSS.n3442 16.0005
R7243 VSS.n3442 VSS.n3441 16.0005
R7244 VSS.n3441 VSS.n3426 16.0005
R7245 VSS.n3427 VSS.n3426 16.0005
R7246 VSS.n3434 VSS.n3427 16.0005
R7247 VSS.n3434 VSS.n3433 16.0005
R7248 VSS.n3433 VSS.n3432 16.0005
R7249 VSS.n3432 VSS.n1274 16.0005
R7250 VSS.n3879 VSS.n1303 16.0005
R7251 VSS.n3880 VSS.n3879 16.0005
R7252 VSS.n3881 VSS.n3880 16.0005
R7253 VSS.n3881 VSS.n1301 16.0005
R7254 VSS.n3886 VSS.n1301 16.0005
R7255 VSS.n3887 VSS.n3886 16.0005
R7256 VSS.n3887 VSS.n1297 16.0005
R7257 VSS.n3892 VSS.n1297 16.0005
R7258 VSS.n4707 VSS.n4704 16.0005
R7259 VSS.n4704 VSS.n4703 16.0005
R7260 VSS.n4703 VSS.n4700 16.0005
R7261 VSS.n4700 VSS.n4699 16.0005
R7262 VSS.n4699 VSS.n4696 16.0005
R7263 VSS.n4696 VSS.n4695 16.0005
R7264 VSS.n4695 VSS.n582 16.0005
R7265 VSS.n5074 VSS.n582 16.0005
R7266 VSS.n722 VSS.n668 16.0005
R7267 VSS.n723 VSS.n722 16.0005
R7268 VSS.n725 VSS.n723 16.0005
R7269 VSS.n726 VSS.n725 16.0005
R7270 VSS.n729 VSS.n726 16.0005
R7271 VSS.n731 VSS.n729 16.0005
R7272 VSS.n732 VSS.n731 16.0005
R7273 VSS.n733 VSS.n732 16.0005
R7274 VSS.n4711 VSS.n4708 16.0005
R7275 VSS.n4712 VSS.n4711 16.0005
R7276 VSS.n4715 VSS.n4712 16.0005
R7277 VSS.n4716 VSS.n4715 16.0005
R7278 VSS.n4719 VSS.n4716 16.0005
R7279 VSS.n4720 VSS.n4719 16.0005
R7280 VSS.n4723 VSS.n4720 16.0005
R7281 VSS.n4773 VSS.n4723 16.0005
R7282 VSS.n4799 VSS.n4796 16.0005
R7283 VSS.n4796 VSS.n4794 16.0005
R7284 VSS.n4794 VSS.n4793 16.0005
R7285 VSS.n4793 VSS.n4791 16.0005
R7286 VSS.n4791 VSS.n4788 16.0005
R7287 VSS.n4788 VSS.n4787 16.0005
R7288 VSS.n4787 VSS.n4785 16.0005
R7289 VSS.n4785 VSS.n4784 16.0005
R7290 VSS.n4819 VSS.n4818 16.0005
R7291 VSS.n4818 VSS.n4817 16.0005
R7292 VSS.n4817 VSS.n665 16.0005
R7293 VSS.n666 VSS.n665 16.0005
R7294 VSS.n4810 VSS.n666 16.0005
R7295 VSS.n4810 VSS.n4809 16.0005
R7296 VSS.n4809 VSS.n4808 16.0005
R7297 VSS.n4808 VSS.n4803 16.0005
R7298 VSS.n4896 VSS.n4895 16.0005
R7299 VSS.n4895 VSS.n4894 16.0005
R7300 VSS.n4894 VSS.n4833 16.0005
R7301 VSS.n4889 VSS.n4833 16.0005
R7302 VSS.n4889 VSS.n4888 16.0005
R7303 VSS.n4888 VSS.n4887 16.0005
R7304 VSS.n4887 VSS.n4836 16.0005
R7305 VSS.n4882 VSS.n4836 16.0005
R7306 VSS.n1843 VSS.n1809 16.0005
R7307 VSS.n1861 VSS.n1843 16.0005
R7308 VSS.n1861 VSS.n1860 16.0005
R7309 VSS.n1860 VSS.n1859 16.0005
R7310 VSS.n1859 VSS.n1845 16.0005
R7311 VSS.n1854 VSS.n1845 16.0005
R7312 VSS.n1854 VSS.n1853 16.0005
R7313 VSS.n1853 VSS.n1852 16.0005
R7314 VSS.n5173 VSS.n5172 16.0005
R7315 VSS.n5172 VSS.n5171 16.0005
R7316 VSS.n5171 VSS.n441 16.0005
R7317 VSS.n5166 VSS.n441 16.0005
R7318 VSS.n5166 VSS.n5165 16.0005
R7319 VSS.n5165 VSS.n5164 16.0005
R7320 VSS.n5164 VSS.n444 16.0005
R7321 VSS.n445 VSS.n444 16.0005
R7322 VSS.n817 VSS.n815 16.0005
R7323 VSS.n818 VSS.n817 16.0005
R7324 VSS.n821 VSS.n818 16.0005
R7325 VSS.n822 VSS.n821 16.0005
R7326 VSS.n825 VSS.n822 16.0005
R7327 VSS.n826 VSS.n825 16.0005
R7328 VSS.n829 VSS.n826 16.0005
R7329 VSS.n830 VSS.n829 16.0005
R7330 VSS.n761 VSS.n758 16.0005
R7331 VSS.n762 VSS.n761 16.0005
R7332 VSS.n765 VSS.n762 16.0005
R7333 VSS.n767 VSS.n765 16.0005
R7334 VSS.n768 VSS.n767 16.0005
R7335 VSS.n770 VSS.n768 16.0005
R7336 VSS.n770 VSS.n769 16.0005
R7337 VSS.n769 VSS.n744 16.0005
R7338 VSS.n4591 VSS.n4589 16.0005
R7339 VSS.n4592 VSS.n4591 16.0005
R7340 VSS.n4594 VSS.n4592 16.0005
R7341 VSS.n4595 VSS.n4594 16.0005
R7342 VSS.n4598 VSS.n4595 16.0005
R7343 VSS.n4600 VSS.n4598 16.0005
R7344 VSS.n4601 VSS.n4600 16.0005
R7345 VSS.n4602 VSS.n4601 16.0005
R7346 VSS.n3176 VSS.n3173 16.0005
R7347 VSS.n3173 VSS.n3172 16.0005
R7348 VSS.n3172 VSS.n3169 16.0005
R7349 VSS.n3169 VSS.n3168 16.0005
R7350 VSS.n3168 VSS.n3166 16.0005
R7351 VSS.n3166 VSS.n3165 16.0005
R7352 VSS.n3165 VSS.n3163 16.0005
R7353 VSS.n3163 VSS.n3160 16.0005
R7354 VSS.n4450 VSS.n4447 16.0005
R7355 VSS.n4451 VSS.n4450 16.0005
R7356 VSS.n4454 VSS.n4451 16.0005
R7357 VSS.n4455 VSS.n4454 16.0005
R7358 VSS.n4458 VSS.n4455 16.0005
R7359 VSS.n4459 VSS.n4458 16.0005
R7360 VSS.n4462 VSS.n4459 16.0005
R7361 VSS.n4505 VSS.n4462 16.0005
R7362 VSS.n4412 VSS.n4410 16.0005
R7363 VSS.n4413 VSS.n4412 16.0005
R7364 VSS.n4415 VSS.n4413 16.0005
R7365 VSS.n4416 VSS.n4415 16.0005
R7366 VSS.n4419 VSS.n4416 16.0005
R7367 VSS.n4421 VSS.n4419 16.0005
R7368 VSS.n4422 VSS.n4421 16.0005
R7369 VSS.n4423 VSS.n4422 16.0005
R7370 VSS.n2363 VSS.n2362 16.0005
R7371 VSS.n2363 VSS.n2065 16.0005
R7372 VSS.n2369 VSS.n2065 16.0005
R7373 VSS.n2370 VSS.n2369 16.0005
R7374 VSS.n2371 VSS.n2370 16.0005
R7375 VSS.n2371 VSS.n2063 16.0005
R7376 VSS.n2376 VSS.n2063 16.0005
R7377 VSS.n2396 VSS.n2376 16.0005
R7378 VSS.n2391 VSS.n2388 16.0005
R7379 VSS.n2388 VSS.n2387 16.0005
R7380 VSS.n2387 VSS.n2384 16.0005
R7381 VSS.n2384 VSS.n2383 16.0005
R7382 VSS.n2383 VSS.n2380 16.0005
R7383 VSS.n2380 VSS.n2379 16.0005
R7384 VSS.n2379 VSS.n2377 16.0005
R7385 VSS.n2377 VSS.n638 16.0005
R7386 VSS.n2031 VSS.n2030 16.0005
R7387 VSS.n2030 VSS.n2028 16.0005
R7388 VSS.n2028 VSS.n2027 16.0005
R7389 VSS.n2027 VSS.n2025 16.0005
R7390 VSS.n2025 VSS.n2022 16.0005
R7391 VSS.n2022 VSS.n2021 16.0005
R7392 VSS.n2021 VSS.n2019 16.0005
R7393 VSS.n2019 VSS.n2018 16.0005
R7394 VSS.n2013 VSS.n2002 16.0005
R7395 VSS.n2443 VSS.n2013 16.0005
R7396 VSS.n2443 VSS.n2442 16.0005
R7397 VSS.n2442 VSS.n2441 16.0005
R7398 VSS.n2441 VSS.n2015 16.0005
R7399 VSS.n2016 VSS.n2015 16.0005
R7400 VSS.n2434 VSS.n2016 16.0005
R7401 VSS.n2434 VSS.n2433 16.0005
R7402 VSS.n2338 VSS.n2113 16.0005
R7403 VSS.n2339 VSS.n2338 16.0005
R7404 VSS.n2340 VSS.n2339 16.0005
R7405 VSS.n2340 VSS.n2111 16.0005
R7406 VSS.n2346 VSS.n2111 16.0005
R7407 VSS.n2347 VSS.n2346 16.0005
R7408 VSS.n2348 VSS.n2347 16.0005
R7409 VSS.n2348 VSS.n2067 16.0005
R7410 VSS.n2151 VSS.n2150 16.0005
R7411 VSS.n2150 VSS.n2132 16.0005
R7412 VSS.n2145 VSS.n2132 16.0005
R7413 VSS.n2145 VSS.n2144 16.0005
R7414 VSS.n2144 VSS.n2134 16.0005
R7415 VSS.n2139 VSS.n2134 16.0005
R7416 VSS.n2139 VSS.n2138 16.0005
R7417 VSS.n2138 VSS.n2003 16.0005
R7418 VSS.n2279 VSS.n2278 16.0005
R7419 VSS.n2278 VSS.n2277 16.0005
R7420 VSS.n2277 VSS.n2255 16.0005
R7421 VSS.n2271 VSS.n2255 16.0005
R7422 VSS.n2271 VSS.n2270 16.0005
R7423 VSS.n2270 VSS.n2269 16.0005
R7424 VSS.n2269 VSS.n2257 16.0005
R7425 VSS.n2257 VSS.n1701 16.0005
R7426 VSS.n2517 VSS.n2516 16.0005
R7427 VSS.n2516 VSS.n1571 16.0005
R7428 VSS.n2512 VSS.n1571 16.0005
R7429 VSS.n2512 VSS.n2511 16.0005
R7430 VSS.n2511 VSS.n1573 16.0005
R7431 VSS.n2506 VSS.n1573 16.0005
R7432 VSS.n2506 VSS.n2505 16.0005
R7433 VSS.n2505 VSS.n2504 16.0005
R7434 VSS.n1556 VSS.n1553 16.0005
R7435 VSS.n1553 VSS.n1552 16.0005
R7436 VSS.n1552 VSS.n1549 16.0005
R7437 VSS.n1549 VSS.n1548 16.0005
R7438 VSS.n1548 VSS.n1545 16.0005
R7439 VSS.n1545 VSS.n1544 16.0005
R7440 VSS.n1544 VSS.n1542 16.0005
R7441 VSS.n1542 VSS.n1456 16.0005
R7442 VSS.n2566 VSS.n2564 16.0005
R7443 VSS.n2567 VSS.n2566 16.0005
R7444 VSS.n2569 VSS.n2567 16.0005
R7445 VSS.n2570 VSS.n2569 16.0005
R7446 VSS.n2573 VSS.n2570 16.0005
R7447 VSS.n2575 VSS.n2573 16.0005
R7448 VSS.n2576 VSS.n2575 16.0005
R7449 VSS.n2577 VSS.n2576 16.0005
R7450 VSS.n5300 VSS.n332 16.0005
R7451 VSS.n5301 VSS.n5300 16.0005
R7452 VSS.n5302 VSS.n5301 16.0005
R7453 VSS.n5302 VSS.n330 16.0005
R7454 VSS.n5308 VSS.n330 16.0005
R7455 VSS.n5309 VSS.n5308 16.0005
R7456 VSS.n5310 VSS.n5309 16.0005
R7457 VSS.n5310 VSS.n328 16.0005
R7458 VSS.n4385 VSS.n4384 16.0005
R7459 VSS.n4384 VSS.n4368 16.0005
R7460 VSS.n4380 VSS.n4368 16.0005
R7461 VSS.n4380 VSS.n4379 16.0005
R7462 VSS.n4379 VSS.n4370 16.0005
R7463 VSS.n4374 VSS.n4370 16.0005
R7464 VSS.n4374 VSS.n4373 16.0005
R7465 VSS.n4373 VSS.n305 16.0005
R7466 VSS.n4183 VSS.n4181 16.0005
R7467 VSS.n4184 VSS.n4183 16.0005
R7468 VSS.n4187 VSS.n4184 16.0005
R7469 VSS.n4188 VSS.n4187 16.0005
R7470 VSS.n4191 VSS.n4188 16.0005
R7471 VSS.n4192 VSS.n4191 16.0005
R7472 VSS.n4195 VSS.n4192 16.0005
R7473 VSS.n4198 VSS.n4195 16.0005
R7474 VSS.n1996 VSS.n1995 16.0005
R7475 VSS.n1995 VSS.n1993 16.0005
R7476 VSS.n1993 VSS.n1990 16.0005
R7477 VSS.n1990 VSS.n1989 16.0005
R7478 VSS.n1989 VSS.n1986 16.0005
R7479 VSS.n1986 VSS.n1985 16.0005
R7480 VSS.n1985 VSS.n1982 16.0005
R7481 VSS.n1982 VSS.n1981 16.0005
R7482 VSS.n1973 VSS.n1972 16.0005
R7483 VSS.n1972 VSS.n1971 16.0005
R7484 VSS.n1971 VSS.n1805 16.0005
R7485 VSS.n1965 VSS.n1805 16.0005
R7486 VSS.n1965 VSS.n1964 16.0005
R7487 VSS.n1964 VSS.n1963 16.0005
R7488 VSS.n1963 VSS.n1807 16.0005
R7489 VSS.n1957 VSS.n1807 16.0005
R7490 VSS.n1762 VSS.n1761 16.0005
R7491 VSS.n1761 VSS.n1743 16.0005
R7492 VSS.n1757 VSS.n1743 16.0005
R7493 VSS.n1757 VSS.n1756 16.0005
R7494 VSS.n1756 VSS.n1745 16.0005
R7495 VSS.n1751 VSS.n1745 16.0005
R7496 VSS.n1751 VSS.n1750 16.0005
R7497 VSS.n1750 VSS.n1749 16.0005
R7498 VSS.n1728 VSS.n1725 16.0005
R7499 VSS.n1729 VSS.n1728 16.0005
R7500 VSS.n1732 VSS.n1729 16.0005
R7501 VSS.n1734 VSS.n1732 16.0005
R7502 VSS.n1735 VSS.n1734 16.0005
R7503 VSS.n1737 VSS.n1735 16.0005
R7504 VSS.n1738 VSS.n1737 16.0005
R7505 VSS.n1741 VSS.n1738 16.0005
R7506 VSS.n3058 VSS.n3057 16.0005
R7507 VSS.n3058 VSS.n1454 16.0005
R7508 VSS.n3064 VSS.n1454 16.0005
R7509 VSS.n3065 VSS.n3064 16.0005
R7510 VSS.n3066 VSS.n3065 16.0005
R7511 VSS.n3066 VSS.n1452 16.0005
R7512 VSS.n3071 VSS.n1452 16.0005
R7513 VSS.n3072 VSS.n3071 16.0005
R7514 VSS.n3092 VSS.n1440 16.0005
R7515 VSS.n3093 VSS.n3092 16.0005
R7516 VSS.n3094 VSS.n3093 16.0005
R7517 VSS.n3094 VSS.n1438 16.0005
R7518 VSS.n3100 VSS.n1438 16.0005
R7519 VSS.n3101 VSS.n3100 16.0005
R7520 VSS.n3102 VSS.n3101 16.0005
R7521 VSS.n3102 VSS.n1436 16.0005
R7522 VSS.n2867 VSS.n2866 16.0005
R7523 VSS.n2866 VSS.n2728 16.0005
R7524 VSS.n2861 VSS.n2728 16.0005
R7525 VSS.n2861 VSS.n2860 16.0005
R7526 VSS.n2860 VSS.n2730 16.0005
R7527 VSS.n2855 VSS.n2730 16.0005
R7528 VSS.n2855 VSS.n2854 16.0005
R7529 VSS.n2854 VSS.n2853 16.0005
R7530 VSS.n2985 VSS.n2984 16.0005
R7531 VSS.n2984 VSS.n2983 16.0005
R7532 VSS.n2983 VSS.n2579 16.0005
R7533 VSS.n2978 VSS.n2579 16.0005
R7534 VSS.n2978 VSS.n2977 16.0005
R7535 VSS.n2977 VSS.n2976 16.0005
R7536 VSS.n2976 VSS.n2582 16.0005
R7537 VSS.n2583 VSS.n2582 16.0005
R7538 VSS.n2704 VSS.n2676 16.0005
R7539 VSS.n2705 VSS.n2704 16.0005
R7540 VSS.n2706 VSS.n2705 16.0005
R7541 VSS.n2706 VSS.n2674 16.0005
R7542 VSS.n2712 VSS.n2674 16.0005
R7543 VSS.n2713 VSS.n2712 16.0005
R7544 VSS.n2714 VSS.n2713 16.0005
R7545 VSS.n2714 VSS.n2622 16.0005
R7546 VSS.n2638 VSS.n2635 16.0005
R7547 VSS.n2635 VSS.n2634 16.0005
R7548 VSS.n2634 VSS.n2631 16.0005
R7549 VSS.n2631 VSS.n2630 16.0005
R7550 VSS.n2630 VSS.n2627 16.0005
R7551 VSS.n2627 VSS.n2626 16.0005
R7552 VSS.n2626 VSS.n2623 16.0005
R7553 VSS.n2623 VSS.n239 16.0005
R7554 VSS.n3269 VSS.n3267 16.0005
R7555 VSS.n3270 VSS.n3269 16.0005
R7556 VSS.n3272 VSS.n3270 16.0005
R7557 VSS.n3273 VSS.n3272 16.0005
R7558 VSS.n3276 VSS.n3273 16.0005
R7559 VSS.n3278 VSS.n3276 16.0005
R7560 VSS.n3279 VSS.n3278 16.0005
R7561 VSS.n3280 VSS.n3279 16.0005
R7562 VSS.n5325 VSS.n306 16.0005
R7563 VSS.n5341 VSS.n5325 16.0005
R7564 VSS.n5341 VSS.n5340 16.0005
R7565 VSS.n5340 VSS.n5339 16.0005
R7566 VSS.n5339 VSS.n5327 16.0005
R7567 VSS.n5328 VSS.n5327 16.0005
R7568 VSS.n5332 VSS.n5328 16.0005
R7569 VSS.n5332 VSS.n5331 16.0005
R7570 VSS.n3127 VSS.n1420 16.0005
R7571 VSS.n3128 VSS.n3127 16.0005
R7572 VSS.n3129 VSS.n3128 16.0005
R7573 VSS.n3129 VSS.n1418 16.0005
R7574 VSS.n3135 VSS.n1418 16.0005
R7575 VSS.n3136 VSS.n3135 16.0005
R7576 VSS.n3137 VSS.n3136 16.0005
R7577 VSS.n3137 VSS.n1389 16.0005
R7578 VSS.n1404 VSS.n1401 16.0005
R7579 VSS.n1401 VSS.n1400 16.0005
R7580 VSS.n1400 VSS.n1397 16.0005
R7581 VSS.n1397 VSS.n1396 16.0005
R7582 VSS.n1396 VSS.n1393 16.0005
R7583 VSS.n1393 VSS.n1392 16.0005
R7584 VSS.n1392 VSS.n1390 16.0005
R7585 VSS.n1390 VSS.n847 16.0005
R7586 VSS.n2787 VSS.n2786 16.0005
R7587 VSS.n2786 VSS.n2784 16.0005
R7588 VSS.n2784 VSS.n2783 16.0005
R7589 VSS.n2783 VSS.n2781 16.0005
R7590 VSS.n2781 VSS.n2778 16.0005
R7591 VSS.n2778 VSS.n2777 16.0005
R7592 VSS.n2777 VSS.n2775 16.0005
R7593 VSS.n2775 VSS.n899 16.0005
R7594 VSS.n2807 VSS.n2806 16.0005
R7595 VSS.n2806 VSS.n2805 16.0005
R7596 VSS.n2805 VSS.n2738 16.0005
R7597 VSS.n2800 VSS.n2738 16.0005
R7598 VSS.n2800 VSS.n2799 16.0005
R7599 VSS.n2799 VSS.n2798 16.0005
R7600 VSS.n2798 VSS.n2741 16.0005
R7601 VSS.n2742 VSS.n2741 16.0005
R7602 VSS.n1326 VSS.n240 16.0005
R7603 VSS.n1327 VSS.n1326 16.0005
R7604 VSS.n1330 VSS.n1327 16.0005
R7605 VSS.n1331 VSS.n1330 16.0005
R7606 VSS.n1334 VSS.n1331 16.0005
R7607 VSS.n1335 VSS.n1334 16.0005
R7608 VSS.n1338 VSS.n1335 16.0005
R7609 VSS.n1341 VSS.n1338 16.0005
R7610 VSS.n3846 VSS.n1322 16.0005
R7611 VSS.n3847 VSS.n3846 16.0005
R7612 VSS.n3848 VSS.n3847 16.0005
R7613 VSS.n3848 VSS.n1320 16.0005
R7614 VSS.n3854 VSS.n1320 16.0005
R7615 VSS.n3855 VSS.n3854 16.0005
R7616 VSS.n3856 VSS.n3855 16.0005
R7617 VSS.n3856 VSS.n1318 16.0005
R7618 VSS.n3492 VSS.n3264 16.0005
R7619 VSS.n3492 VSS.n3491 16.0005
R7620 VSS.n3491 VSS.n3490 16.0005
R7621 VSS.n3490 VSS.n3415 16.0005
R7622 VSS.n3485 VSS.n3415 16.0005
R7623 VSS.n3485 VSS.n3484 16.0005
R7624 VSS.n3484 VSS.n3417 16.0005
R7625 VSS.n3418 VSS.n3417 16.0005
R7626 VSS.n3353 VSS.n3350 16.0005
R7627 VSS.n3354 VSS.n3353 16.0005
R7628 VSS.n3357 VSS.n3354 16.0005
R7629 VSS.n3359 VSS.n3357 16.0005
R7630 VSS.n3360 VSS.n3359 16.0005
R7631 VSS.n3362 VSS.n3360 16.0005
R7632 VSS.n3363 VSS.n3362 16.0005
R7633 VSS.n3366 VSS.n3363 16.0005
R7634 VSS.n4043 VSS.n4040 16.0005
R7635 VSS.n4040 VSS.n4037 16.0005
R7636 VSS.n4037 VSS.n4036 16.0005
R7637 VSS.n4036 VSS.n4033 16.0005
R7638 VSS.n4033 VSS.n4032 16.0005
R7639 VSS.n4032 VSS.n4029 16.0005
R7640 VSS.n4029 VSS.n4028 16.0005
R7641 VSS.n4028 VSS.n4025 16.0005
R7642 VSS.n4063 VSS.n1108 16.0005
R7643 VSS.n4057 VSS.n1108 16.0005
R7644 VSS.n4057 VSS.n4056 16.0005
R7645 VSS.n4056 VSS.n4055 16.0005
R7646 VSS.n4055 VSS.n1110 16.0005
R7647 VSS.n1111 VSS.n1110 16.0005
R7648 VSS.n4048 VSS.n1111 16.0005
R7649 VSS.n4048 VSS.n4047 16.0005
R7650 VSS.n4122 VSS.n4121 16.0005
R7651 VSS.n4125 VSS.n4122 16.0005
R7652 VSS.n4126 VSS.n4125 16.0005
R7653 VSS.n4129 VSS.n4126 16.0005
R7654 VSS.n4130 VSS.n4129 16.0005
R7655 VSS.n4133 VSS.n4130 16.0005
R7656 VSS.n4134 VSS.n4133 16.0005
R7657 VSS.n4137 VSS.n4134 16.0005
R7658 VSS.n4107 VSS.n4105 16.0005
R7659 VSS.n4108 VSS.n4107 16.0005
R7660 VSS.n4110 VSS.n4108 16.0005
R7661 VSS.n4111 VSS.n4110 16.0005
R7662 VSS.n4114 VSS.n4111 16.0005
R7663 VSS.n4116 VSS.n4114 16.0005
R7664 VSS.n4117 VSS.n4116 16.0005
R7665 VSS.n4118 VSS.n4117 16.0005
R7666 VSS.n3998 VSS.n3997 15.5797
R7667 VSS.n5286 VSS.n342 15.0432
R7668 VSS.n5567 VSS.n0 14.6031
R7669 VSS.n3800 VSS.n3522 13.6894
R7670 VSS.n3705 VSS.n3704 13.6894
R7671 VSS.n1303 VSS.n901 13.6894
R7672 VSS.n4775 VSS.n4707 13.6894
R7673 VSS.n815 VSS.n485 13.6894
R7674 VSS.n758 VSS.n669 13.6894
R7675 VSS.n4447 VSS.n4446 13.6894
R7676 VSS.n3159 VSS.n1404 13.6894
R7677 VSS.n1342 VSS.n1322 13.6894
R7678 VSS.n25 VSS.n15 13.6602
R7679 VSS.n2117 VSS.n2113 13.5116
R7680 VSS.n2279 VSS.n2222 13.5116
R7681 VSS.n1557 VSS.n1556 13.5116
R7682 VSS.n335 VSS.n332 13.5116
R7683 VSS.n4181 VSS.n1013 13.5116
R7684 VSS.n1145 VSS.t101 13.3541
R7685 VSS.n4199 VSS.n4180 13.3338
R7686 VSS.n5430 VSS.n5429 13.3338
R7687 VSS.n3507 VSS.n113 13.3338
R7688 VSS.n4896 VSS.n4832 13.3338
R7689 VSS.n1956 VSS.n1809 13.3338
R7690 VSS.n2362 VSS.n2361 13.3338
R7691 VSS.n2395 VSS.n2391 13.3338
R7692 VSS.n2470 VSS.n1996 13.3338
R7693 VSS.n1973 VSS.n1702 13.3338
R7694 VSS.n3057 VSS.n3056 13.3338
R7695 VSS.n1443 VSS.n1440 13.3338
R7696 VSS.n2676 VSS.n295 13.3338
R7697 VSS.n2727 VSS.n2638 13.3338
R7698 VSS.n1435 VSS.n1420 13.3338
R7699 VSS.n5377 VSS.n240 13.3338
R7700 VSS.n4708 VSS.n607 13.1561
R7701 VSS.n5493 VSS.t25 11.6849
R7702 VSS.n5479 VSS.t3 11.6849
R7703 VSS.n11 VSS.n9 11.6369
R7704 VSS.n5554 VSS.n11 11.6369
R7705 VSS.n5554 VSS.n5553 11.6369
R7706 VSS.n5553 VSS.n5552 11.6369
R7707 VSS.n5552 VSS.n12 11.6369
R7708 VSS.n5546 VSS.n12 11.6369
R7709 VSS.n5546 VSS.n5545 11.6369
R7710 VSS.n5545 VSS.n5544 11.6369
R7711 VSS.n5497 VSS.n62 11.6369
R7712 VSS.n5491 VSS.n62 11.6369
R7713 VSS.n5491 VSS.n5490 11.6369
R7714 VSS.n5490 VSS.n5489 11.6369
R7715 VSS.n5489 VSS.n66 11.6369
R7716 VSS.n5483 VSS.n66 11.6369
R7717 VSS.n5483 VSS.n5482 11.6369
R7718 VSS.n5482 VSS.n5481 11.6369
R7719 VSS.n5532 VSS.n5531 11.6369
R7720 VSS.n5531 VSS.n5530 11.6369
R7721 VSS.n5530 VSS.n36 11.6369
R7722 VSS.n5524 VSS.n36 11.6369
R7723 VSS.n5524 VSS.n5523 11.6369
R7724 VSS.n5523 VSS.n5522 11.6369
R7725 VSS.n5522 VSS.n41 11.6369
R7726 VSS.n5516 VSS.n41 11.6369
R7727 VSS.n4003 VSS.n4002 11.6369
R7728 VSS.n4002 VSS.n4001 11.6369
R7729 VSS.n4001 VSS.n1197 11.6369
R7730 VSS.n1206 VSS.n1197 11.6369
R7731 VSS.n1208 VSS.n1206 11.6369
R7732 VSS.n1208 VSS.n1207 11.6369
R7733 VSS.n1207 VSS.n1203 11.6369
R7734 VSS.n1215 VSS.n1203 11.6369
R7735 VSS.n4997 VSS.n624 11.6369
R7736 VSS.n4998 VSS.n4997 11.6369
R7737 VSS.n4999 VSS.n4998 11.6369
R7738 VSS.n4999 VSS.n618 11.6369
R7739 VSS.n5005 VSS.n618 11.6369
R7740 VSS.n5006 VSS.n5005 11.6369
R7741 VSS.n5007 VSS.n5006 11.6369
R7742 VSS.n5007 VSS.n608 11.6369
R7743 VSS.n355 VSS.n352 11.6369
R7744 VSS.n5272 VSS.n355 11.6369
R7745 VSS.n5272 VSS.n5271 11.6369
R7746 VSS.n5271 VSS.n5270 11.6369
R7747 VSS.n5270 VSS.n356 11.6369
R7748 VSS.n5264 VSS.n356 11.6369
R7749 VSS.n5264 VSS.n5263 11.6369
R7750 VSS.n5263 VSS.n5262 11.6369
R7751 VSS.n4970 VSS.n4968 11.6369
R7752 VSS.n4970 VSS.n4969 11.6369
R7753 VSS.n4969 VSS.n4959 11.6369
R7754 VSS.n4959 VSS.n4957 11.6369
R7755 VSS.n4980 VSS.n4957 11.6369
R7756 VSS.n4981 VSS.n4980 11.6369
R7757 VSS.n4983 VSS.n4981 11.6369
R7758 VSS.n4983 VSS.n4982 11.6369
R7759 VSS.n5249 VSS.n370 11.6369
R7760 VSS.n5249 VSS.n5248 11.6369
R7761 VSS.n5248 VSS.n5247 11.6369
R7762 VSS.n5247 VSS.n371 11.6369
R7763 VSS.n5241 VSS.n371 11.6369
R7764 VSS.n5241 VSS.n5240 11.6369
R7765 VSS.n5240 VSS.n5239 11.6369
R7766 VSS.n5239 VSS.n377 11.6369
R7767 VSS.n5017 VSS.n603 11.6369
R7768 VSS.n5024 VSS.n603 11.6369
R7769 VSS.n5025 VSS.n5024 11.6369
R7770 VSS.n5026 VSS.n5025 11.6369
R7771 VSS.n5026 VSS.n600 11.6369
R7772 VSS.n5032 VSS.n600 11.6369
R7773 VSS.n5033 VSS.n5032 11.6369
R7774 VSS.n5035 VSS.n5033 11.6369
R7775 VSS.n5035 VSS.n5034 11.6369
R7776 VSS.n5034 VSS.n597 11.6369
R7777 VSS.n5045 VSS.n5044 11.6369
R7778 VSS.n5046 VSS.n5045 11.6369
R7779 VSS.n5046 VSS.n590 11.6369
R7780 VSS.n5053 VSS.n590 11.6369
R7781 VSS.n5054 VSS.n5053 11.6369
R7782 VSS.n5055 VSS.n5054 11.6369
R7783 VSS.n5055 VSS.n587 11.6369
R7784 VSS.n5062 VSS.n587 11.6369
R7785 VSS.n5063 VSS.n5062 11.6369
R7786 VSS.n5064 VSS.n5063 11.6369
R7787 VSS.n1141 VSS.n1132 11.6369
R7788 VSS.n1142 VSS.n1141 11.6369
R7789 VSS.n1158 VSS.n1142 11.6369
R7790 VSS.n1158 VSS.n1157 11.6369
R7791 VSS.n1157 VSS.n1156 11.6369
R7792 VSS.n1156 VSS.n1143 11.6369
R7793 VSS.n1150 VSS.n1143 11.6369
R7794 VSS.n1150 VSS.n1149 11.6369
R7795 VSS.n3729 VSS.n3720 11.6369
R7796 VSS.n3730 VSS.n3729 11.6369
R7797 VSS.n3731 VSS.n3730 11.6369
R7798 VSS.n3731 VSS.n3716 11.6369
R7799 VSS.n3738 VSS.n3716 11.6369
R7800 VSS.n3739 VSS.n3738 11.6369
R7801 VSS.n3741 VSS.n3739 11.6369
R7802 VSS.n3741 VSS.n3740 11.6369
R7803 VSS.n3740 VSS.n3713 11.6369
R7804 VSS.n2928 VSS.n2927 11.5043
R7805 VSS.n945 VSS.n902 11.5043
R7806 VSS.n2816 VSS.n2815 11.5043
R7807 VSS.n2995 VSS.n2994 11.5043
R7808 VSS.n4003 VSS.n1196 11.0106
R7809 VSS.n5498 VSS.n5497 10.9261
R7810 VSS.n3748 VSS.n3713 10.9063
R7811 VSS.n4968 VSS.n4967 10.8998
R7812 VSS.t93 VSS.n38 10.5721
R7813 VSS.n4024 VSS.n1114 10.3116
R7814 VSS.n3761 VSS.n3578 10.3116
R7815 VSS.n3443 VSS.n3425 10.3116
R7816 VSS.n4783 VSS.n668 10.3116
R7817 VSS.n4802 VSS.n4799 10.3116
R7818 VSS.n4589 VSS.n786 10.3116
R7819 VSS.n3177 VSS.n3176 10.3116
R7820 VSS.n4410 VSS.n4409 10.3116
R7821 VSS.n2787 VSS.n2774 10.3116
R7822 VSS.n3506 VSS.n3264 10.3116
R7823 VSS.n2152 VSS.n2151 10.1338
R7824 VSS.n2517 VSS.n1562 10.1338
R7825 VSS.n2564 VSS.n1488 10.1338
R7826 VSS.n4385 VSS.n4332 10.1338
R7827 VSS.n4105 VSS.n4066 10.1338
R7828 VSS.n352 VSS.n350 10.0645
R7829 VSS.t14 VSS.n5557 10.0157
R7830 VSS.n1139 VSS.t16 10.0157
R7831 VSS.n9 VSS.n7 9.95606
R7832 VSS.n4819 VSS.n664 9.95606
R7833 VSS.n5173 VSS.n440 9.95606
R7834 VSS.n2432 VSS.n2031 9.95606
R7835 VSS.n2464 VSS.n2002 9.95606
R7836 VSS.n1762 VSS.n1742 9.95606
R7837 VSS.n1725 VSS.n1575 9.95606
R7838 VSS.n2868 VSS.n2867 9.95606
R7839 VSS.n2985 VSS.n2578 9.95606
R7840 VSS.n3267 VSS.n148 9.95606
R7841 VSS.n5361 VSS.n306 9.95606
R7842 VSS.n2807 VSS.n2733 9.95606
R7843 VSS.n3350 VSS.n3349 9.95606
R7844 VSS.n4046 VSS.n4043 9.95606
R7845 VSS.n4138 VSS.n4063 9.95606
R7846 VSS.n4121 VSS.n4120 9.95606
R7847 VSS.n5532 VSS.n28 9.82676
R7848 VSS.n4952 VSS.n624 9.82676
R7849 VSS.n370 VSS.n360 9.82676
R7850 VSS.n5017 VSS.n5016 9.82676
R7851 VSS.n1132 VSS.n71 9.82676
R7852 VSS.n3723 VSS.n3720 9.80931
R7853 VSS.n597 VSS.n594 9.69747
R7854 VSS.n1139 VSS.t31 9.45928
R7855 VSS.n3988 VSS.n1219 8.95269
R7856 VSS.n1147 VSS.t23 8.90288
R7857 VSS.n18 VSS.t15 8.7005
R7858 VSS.n18 VSS.t66 8.7005
R7859 VSS.n16 VSS.t11 8.7005
R7860 VSS.n16 VSS.t13 8.7005
R7861 VSS.n5516 VSS.n5515 8.13406
R7862 VSS.n1149 VSS.n1127 8.08329
R7863 VSS.n5233 VSS.n377 8.00427
R7864 VSS.n3762 VSS.n3761 7.11161
R7865 VSS.n3991 VSS.n1216 7.11161
R7866 VSS.n3955 VSS.n1274 7.11161
R7867 VSS.n734 VSS.n733 7.11161
R7868 VSS.n4784 VSS.n4783 7.11161
R7869 VSS.n4803 VSS.n4802 7.11161
R7870 VSS.n3177 VSS.n445 7.11161
R7871 VSS.n4603 VSS.n4602 7.11161
R7872 VSS.n3160 VSS.n786 7.11161
R7873 VSS.n4424 VSS.n4423 7.11161
R7874 VSS.n2433 VSS.n2432 7.11161
R7875 VSS.n1742 VSS.n1741 7.11161
R7876 VSS.n2868 VSS.n2583 7.11161
R7877 VSS.n5331 VSS.n148 7.11161
R7878 VSS.n4409 VSS.n899 7.11161
R7879 VSS.n2774 VSS.n2742 7.11161
R7880 VSS.n3425 VSS.n3418 7.11161
R7881 VSS.n3506 VSS.n3366 7.11161
R7882 VSS.n4025 VSS.n4024 7.11161
R7883 VSS.n4138 VSS.n4137 7.11161
R7884 VSS.n5515 VSS.n5514 7.06798
R7885 VSS.n5499 VSS.n5498 7.06798
R7886 VSS.n4017 VSS.n1127 7.06798
R7887 VSS.n3749 VSS.n3748 6.94026
R7888 VSS.n3755 VSS.n1196 6.94026
R7889 VSS.n2018 VSS.n664 6.93383
R7890 VSS.n2464 VSS.n2003 6.93383
R7891 VSS.n2504 VSS.n1575 6.93383
R7892 VSS.n2578 VSS.n2577 6.93383
R7893 VSS.n5361 VSS.n305 6.93383
R7894 VSS.n1749 VSS.n440 6.93383
R7895 VSS.n2853 VSS.n2733 6.93383
R7896 VSS.n3349 VSS.n3280 6.93383
R7897 VSS.n4047 VSS.n4046 6.93383
R7898 VSS.n4120 VSS.n4118 6.93383
R7899 VSS.n5233 VSS.n5232 6.8987
R7900 VSS.n4967 VSS.n4962 6.8987
R7901 VSS.n5499 VSS.n61 6.59682
R7902 VSS.n3723 VSS.n1126 6.59682
R7903 VSS.n3756 VSS.n3755 6.47761
R7904 VSS.n1126 VSS.n1115 6.43976
R7905 VSS.n4962 VSS.n383 6.43882
R7906 VSS.n3711 VSS.n3579 6.16917
R7907 VSS.n1249 VSS.n1245 5.81868
R7908 VSS.n1250 VSS.n1249 5.81868
R7909 VSS.n1254 VSS.n1250 5.81868
R7910 VSS.n1255 VSS.n1254 5.81868
R7911 VSS.n1259 VSS.n1255 5.81868
R7912 VSS.n1260 VSS.n1259 5.81868
R7913 VSS.n1264 VSS.n1260 5.81868
R7914 VSS.n1267 VSS.n1264 5.81868
R7915 VSS.n4478 VSS.n4469 5.81868
R7916 VSS.n4479 VSS.n4478 5.81868
R7917 VSS.n4479 VSS.n4467 5.81868
R7918 VSS.n4485 VSS.n4467 5.81868
R7919 VSS.n4486 VSS.n4485 5.81868
R7920 VSS.n4486 VSS.n4465 5.81868
R7921 VSS.n4492 VSS.n4465 5.81868
R7922 VSS.n4494 VSS.n4492 5.81868
R7923 VSS.n3180 VSS.n3179 5.81868
R7924 VSS.n3208 VSS.n3180 5.81868
R7925 VSS.n3208 VSS.n3207 5.81868
R7926 VSS.n3207 VSS.n3182 5.81868
R7927 VSS.n3183 VSS.n3182 5.81868
R7928 VSS.n3199 VSS.n3183 5.81868
R7929 VSS.n3199 VSS.n3198 5.81868
R7930 VSS.n3198 VSS.n3185 5.81868
R7931 VSS.n3186 VSS.n3185 5.81868
R7932 VSS.n3902 VSS.n3901 5.81868
R7933 VSS.n3906 VSS.n3902 5.81868
R7934 VSS.n3907 VSS.n3906 5.81868
R7935 VSS.n3911 VSS.n3907 5.81868
R7936 VSS.n3912 VSS.n3911 5.81868
R7937 VSS.n3916 VSS.n3912 5.81868
R7938 VSS.n3917 VSS.n3916 5.81868
R7939 VSS.n3921 VSS.n3917 5.81868
R7940 VSS.n2896 VSS.n2893 5.81868
R7941 VSS.n2893 VSS.n2889 5.81868
R7942 VSS.n2889 VSS.n2888 5.81868
R7943 VSS.n2888 VSS.n2884 5.81868
R7944 VSS.n2884 VSS.n2883 5.81868
R7945 VSS.n2883 VSS.n2879 5.81868
R7946 VSS.n2879 VSS.n2878 5.81868
R7947 VSS.n2878 VSS.n2874 5.81868
R7948 VSS.n2198 VSS.n2164 5.81868
R7949 VSS.n2168 VSS.n2164 5.81868
R7950 VSS.n2190 VSS.n2168 5.81868
R7951 VSS.n2190 VSS.n2189 5.81868
R7952 VSS.n2189 VSS.n2170 5.81868
R7953 VSS.n2171 VSS.n2170 5.81868
R7954 VSS.n2181 VSS.n2171 5.81868
R7955 VSS.n2181 VSS.n2180 5.81868
R7956 VSS.n1932 VSS.n1931 5.81868
R7957 VSS.n1932 VSS.n1923 5.81868
R7958 VSS.n1938 VSS.n1923 5.81868
R7959 VSS.n1939 VSS.n1938 5.81868
R7960 VSS.n1939 VSS.n1921 5.81868
R7961 VSS.n1945 VSS.n1921 5.81868
R7962 VSS.n1946 VSS.n1945 5.81868
R7963 VSS.n1946 VSS.n1880 5.81868
R7964 VSS.n1910 VSS.n1881 5.81868
R7965 VSS.n1910 VSS.n1909 5.81868
R7966 VSS.n1909 VSS.n1884 5.81868
R7967 VSS.n1885 VSS.n1884 5.81868
R7968 VSS.n1901 VSS.n1885 5.81868
R7969 VSS.n1901 VSS.n1900 5.81868
R7970 VSS.n1900 VSS.n1887 5.81868
R7971 VSS.n1888 VSS.n1887 5.81868
R7972 VSS.n4678 VSS.n712 5.81868
R7973 VSS.n713 VSS.n712 5.81868
R7974 VSS.n4670 VSS.n713 5.81868
R7975 VSS.n4670 VSS.n4669 5.81868
R7976 VSS.n4669 VSS.n715 5.81868
R7977 VSS.n716 VSS.n715 5.81868
R7978 VSS.n4661 VSS.n716 5.81868
R7979 VSS.n4661 VSS.n4660 5.81868
R7980 VSS.n2216 VSS.n2155 5.81868
R7981 VSS.n2216 VSS.n2215 5.81868
R7982 VSS.n2215 VSS.n2157 5.81868
R7983 VSS.n2158 VSS.n2157 5.81868
R7984 VSS.n2207 VSS.n2158 5.81868
R7985 VSS.n2207 VSS.n2206 5.81868
R7986 VSS.n2206 VSS.n2160 5.81868
R7987 VSS.n2200 VSS.n2160 5.81868
R7988 VSS.n1661 VSS.n1560 5.81868
R7989 VSS.n1662 VSS.n1661 5.81868
R7990 VSS.n1662 VSS.n1655 5.81868
R7991 VSS.n1668 VSS.n1655 5.81868
R7992 VSS.n1669 VSS.n1668 5.81868
R7993 VSS.n1669 VSS.n1653 5.81868
R7994 VSS.n1675 VSS.n1653 5.81868
R7995 VSS.n1676 VSS.n1675 5.81868
R7996 VSS.n1516 VSS.n1513 5.81868
R7997 VSS.n1513 VSS.n1509 5.81868
R7998 VSS.n1509 VSS.n1508 5.81868
R7999 VSS.n1508 VSS.n1504 5.81868
R8000 VSS.n1504 VSS.n1503 5.81868
R8001 VSS.n1503 VSS.n1499 5.81868
R8002 VSS.n1499 VSS.n1498 5.81868
R8003 VSS.n1498 VSS.n1494 5.81868
R8004 VSS.n4205 VSS.n1012 5.81868
R8005 VSS.n4209 VSS.n4205 5.81868
R8006 VSS.n4210 VSS.n4209 5.81868
R8007 VSS.n4214 VSS.n4210 5.81868
R8008 VSS.n4215 VSS.n4214 5.81868
R8009 VSS.n4219 VSS.n4215 5.81868
R8010 VSS.n4220 VSS.n4219 5.81868
R8011 VSS.n4224 VSS.n4220 5.81868
R8012 VSS.n2918 VSS.n2917 5.81868
R8013 VSS.n2917 VSS.n2913 5.81868
R8014 VSS.n2913 VSS.n2912 5.81868
R8015 VSS.n2912 VSS.n2908 5.81868
R8016 VSS.n2908 VSS.n2907 5.81868
R8017 VSS.n2907 VSS.n2903 5.81868
R8018 VSS.n2903 VSS.n2902 5.81868
R8019 VSS.n2902 VSS.n2898 5.81868
R8020 VSS.n2597 VSS.n2596 5.81868
R8021 VSS.n2601 VSS.n2597 5.81868
R8022 VSS.n2602 VSS.n2601 5.81868
R8023 VSS.n2606 VSS.n2602 5.81868
R8024 VSS.n2607 VSS.n2606 5.81868
R8025 VSS.n2611 VSS.n2607 5.81868
R8026 VSS.n2612 VSS.n2611 5.81868
R8027 VSS.n2616 VSS.n2612 5.81868
R8028 VSS.n5214 VSS.n408 5.81868
R8029 VSS.n5214 VSS.n5213 5.81868
R8030 VSS.n5213 VSS.n410 5.81868
R8031 VSS.n411 VSS.n410 5.81868
R8032 VSS.n5205 VSS.n411 5.81868
R8033 VSS.n5205 VSS.n5204 5.81868
R8034 VSS.n5204 VSS.n413 5.81868
R8035 VSS.n5198 VSS.n413 5.81868
R8036 VSS.n1643 VSS.n1615 5.81868
R8037 VSS.n1643 VSS.n1642 5.81868
R8038 VSS.n1642 VSS.n1617 5.81868
R8039 VSS.n1618 VSS.n1617 5.81868
R8040 VSS.n1634 VSS.n1618 5.81868
R8041 VSS.n1634 VSS.n1633 5.81868
R8042 VSS.n1633 VSS.n1620 5.81868
R8043 VSS.n1621 VSS.n1620 5.81868
R8044 VSS.n3253 VSS.n3249 5.81868
R8045 VSS.n3249 VSS.n3248 5.81868
R8046 VSS.n3248 VSS.n3244 5.81868
R8047 VSS.n3244 VSS.n3243 5.81868
R8048 VSS.n3243 VSS.n3239 5.81868
R8049 VSS.n3239 VSS.n3238 5.81868
R8050 VSS.n3238 VSS.n3234 5.81868
R8051 VSS.n3234 VSS.n3233 5.81868
R8052 VSS.n3233 VSS.n3229 5.81868
R8053 VSS.n1365 VSS.n415 5.81868
R8054 VSS.n1365 VSS.n1361 5.81868
R8055 VSS.n1371 VSS.n1361 5.81868
R8056 VSS.n1372 VSS.n1371 5.81868
R8057 VSS.n1372 VSS.n1359 5.81868
R8058 VSS.n1378 VSS.n1359 5.81868
R8059 VSS.n1379 VSS.n1378 5.81868
R8060 VSS.n1379 VSS.n1357 5.81868
R8061 VSS.n687 VSS.n685 5.81868
R8062 VSS.n688 VSS.n687 5.81868
R8063 VSS.n692 VSS.n688 5.81868
R8064 VSS.n693 VSS.n692 5.81868
R8065 VSS.n697 VSS.n693 5.81868
R8066 VSS.n698 VSS.n697 5.81868
R8067 VSS.n702 VSS.n698 5.81868
R8068 VSS.n704 VSS.n702 5.81868
R8069 VSS.n707 VSS.n704 5.81868
R8070 VSS.n3830 VSS.n3826 5.81868
R8071 VSS.n3826 VSS.n3825 5.81868
R8072 VSS.n3825 VSS.n3821 5.81868
R8073 VSS.n3821 VSS.n3820 5.81868
R8074 VSS.n3820 VSS.n3816 5.81868
R8075 VSS.n3816 VSS.n3815 5.81868
R8076 VSS.n3815 VSS.n3811 5.81868
R8077 VSS.n3811 VSS.n3810 5.81868
R8078 VSS.n3810 VSS.n3806 5.81868
R8079 VSS.n3307 VSS.n3303 5.81868
R8080 VSS.n3303 VSS.n3302 5.81868
R8081 VSS.n3302 VSS.n3298 5.81868
R8082 VSS.n3298 VSS.n3297 5.81868
R8083 VSS.n3297 VSS.n3293 5.81868
R8084 VSS.n3293 VSS.n3292 5.81868
R8085 VSS.n3292 VSS.n3288 5.81868
R8086 VSS.n3288 VSS.n3287 5.81868
R8087 VSS.n3313 VSS.n3312 5.81868
R8088 VSS.n3317 VSS.n3313 5.81868
R8089 VSS.n3318 VSS.n3317 5.81868
R8090 VSS.n3322 VSS.n3318 5.81868
R8091 VSS.n3323 VSS.n3322 5.81868
R8092 VSS.n3327 VSS.n3323 5.81868
R8093 VSS.n3328 VSS.n3327 5.81868
R8094 VSS.n3332 VSS.n3328 5.81868
R8095 VSS.n4251 VSS.n4247 5.81868
R8096 VSS.n4247 VSS.n4246 5.81868
R8097 VSS.n4246 VSS.n4242 5.81868
R8098 VSS.n4242 VSS.n4241 5.81868
R8099 VSS.n4241 VSS.n4237 5.81868
R8100 VSS.n4237 VSS.n4236 5.81868
R8101 VSS.n4236 VSS.n4232 5.81868
R8102 VSS.n4232 VSS.n4231 5.81868
R8103 VSS.t42 VSS.n1124 5.56449
R8104 VSS.n1245 VSS.n961 5.51409
R8105 VSS.n4472 VSS.n4469 5.51409
R8106 VSS.n3901 VSS.n3897 5.51409
R8107 VSS.n4679 VSS.n4678 5.51409
R8108 VSS.n3993 VSS.n3992 5.50178
R8109 VSS.n3956 VSS.n1271 5.50178
R8110 VSS.n4425 VSS.n898 5.50178
R8111 VSS.n4604 VSS.n785 5.50178
R8112 VSS.n4656 VSS.n4655 5.50178
R8113 VSS.n57 VSS.n56 5.48621
R8114 VSS.n4065 VSS.n7 5.47847
R8115 VSS.n4398 VSS.n4397 5.47847
R8116 VSS.n1522 VSS.n1521 5.47847
R8117 VSS.n2531 VSS.n2529 5.47847
R8118 VSS.n2295 VSS.n2294 5.47847
R8119 VSS.n3190 VSS.n3186 5.46332
R8120 VSS.n1931 VSS.n1925 5.46332
R8121 VSS.n2922 VSS.n2918 5.46332
R8122 VSS.n408 VSS.n405 5.46332
R8123 VSS.n3229 VSS.n3228 5.46332
R8124 VSS.n707 VSS.n706 5.46332
R8125 VSS.n3806 VSS.n3805 5.46332
R8126 VSS.n3312 VSS.n3308 5.46332
R8127 VSS.n1165 VSS.n1163 5.27109
R8128 VSS.n1269 VSS.n1268 5.22944
R8129 VSS.n3924 VSS.n3923 5.22944
R8130 VSS.n4503 VSS.n4463 5.22944
R8131 VSS.n737 VSS.n736 5.22944
R8132 VSS.n5072 VSS.n583 5.22944
R8133 VSS.n4330 VSS.n4329 5.20728
R8134 VSS.n1519 VSS.n1517 5.20728
R8135 VSS.n2534 VSS.n2533 5.20728
R8136 VSS.n2291 VSS.n2290 5.20728
R8137 VSS.n2116 VSS.n350 5.20728
R8138 VSS.n2155 VSS.n2154 4.97828
R8139 VSS.n2532 VSS.n1560 4.97828
R8140 VSS.n1520 VSS.n1516 4.97828
R8141 VSS.n4331 VSS.n1012 4.97828
R8142 VSS.n2897 VSS.n2896 4.91363
R8143 VSS.n2199 VSS.n2198 4.91363
R8144 VSS.n1953 VSS.n1881 4.91363
R8145 VSS.n2596 VSS.n293 4.91363
R8146 VSS.n1615 VSS.n1613 4.91363
R8147 VSS.n5197 VSS.n415 4.91363
R8148 VSS.n3333 VSS.n3307 4.91363
R8149 VSS.n4252 VSS.n4251 4.91363
R8150 VSS.n3216 VSS.n3179 4.90491
R8151 VSS.n3255 VSS.n3253 4.90491
R8152 VSS.n685 VSS.n501 4.90491
R8153 VSS.n3832 VSS.n3830 4.90491
R8154 VSS.n59 VSS.t17 4.45169
R8155 VSS.n1161 VSS.n1129 4.45169
R8156 VSS.n4012 VSS.n4011 4.32991
R8157 VSS.n4064 VSS.n45 4.24099
R8158 VSS.n2394 VSS.n381 4.13942
R8159 VSS.n2180 VSS.n2173 4.06728
R8160 VSS.n2619 VSS.n2616 4.06728
R8161 VSS.n1625 VSS.n1621 4.06728
R8162 VSS.n4231 VSS.n4227 4.06728
R8163 VSS.n2874 VSS.n2873 4.0419
R8164 VSS.n1892 VSS.n1888 4.0419
R8165 VSS.n1385 VSS.n1357 4.0419
R8166 VSS.n3287 VSS.n3283 4.0419
R8167 VSS.n1222 VSS.n1217 4.03114
R8168 VSS.n3984 VSS.n1223 4.03114
R8169 VSS.n3983 VSS.n1224 4.03114
R8170 VSS.n1228 VSS.n1226 4.03114
R8171 VSS.n3978 VSS.n3977 4.03114
R8172 VSS.n3971 VSS.n1236 4.03114
R8173 VSS.n3970 VSS.n1237 4.03114
R8174 VSS.n3966 VSS.n3965 4.03114
R8175 VSS.n3953 VSS.n1275 4.03114
R8176 VSS.n1279 VSS.n1277 4.03114
R8177 VSS.n3948 VSS.n3947 4.03114
R8178 VSS.n3939 VSS.n1280 4.03114
R8179 VSS.n3938 VSS.n1283 4.03114
R8180 VSS.n3933 VSS.n3932 4.03114
R8181 VSS.n1295 VSS.n1288 4.03114
R8182 VSS.n3926 VSS.n1296 4.03114
R8183 VSS.n4531 VSS.n4530 4.03114
R8184 VSS.n4431 VSS.n893 4.03114
R8185 VSS.n4524 VSS.n4432 4.03114
R8186 VSS.n4523 VSS.n4520 4.03114
R8187 VSS.n4519 VSS.n4433 4.03114
R8188 VSS.n4440 VSS.n4434 4.03114
R8189 VSS.n4509 VSS.n4443 4.03114
R8190 VSS.n4508 VSS.n4444 4.03114
R8191 VSS.n4637 VSS.n4636 4.03114
R8192 VSS.n4610 VSS.n780 4.03114
R8193 VSS.n4630 VSS.n4611 4.03114
R8194 VSS.n4629 VSS.n4626 4.03114
R8195 VSS.n4625 VSS.n4612 4.03114
R8196 VSS.n4616 VSS.n4613 4.03114
R8197 VSS.n4644 VSS.n740 4.03114
R8198 VSS.n4643 VSS.n741 4.03114
R8199 VSS.n5100 VSS.n5099 4.03114
R8200 VSS.n568 VSS.n562 4.03114
R8201 VSS.n5093 VSS.n569 4.03114
R8202 VSS.n5092 VSS.n5089 4.03114
R8203 VSS.n5088 VSS.n570 4.03114
R8204 VSS.n577 VSS.n571 4.03114
R8205 VSS.n5078 VSS.n580 4.03114
R8206 VSS.n5077 VSS.n581 4.03114
R8207 VSS.n5487 VSS.t44 3.89529
R8208 VSS.n5508 VSS.n5507 3.77317
R8209 VSS.n5429 VSS.n146 3.73383
R8210 VSS.n3800 VSS.n3521 3.73383
R8211 VSS.n3705 VSS.n3608 3.73383
R8212 VSS.n3690 VSS.n1241 3.73383
R8213 VSS.n3925 VSS.n3892 3.73383
R8214 VSS.n5074 VSS.n5073 3.73383
R8215 VSS.n4775 VSS.n4773 3.73383
R8216 VSS.n4882 VSS.n4881 3.73383
R8217 VSS.n1852 VSS.n485 3.73383
R8218 VSS.n830 VSS.n669 3.73383
R8219 VSS.n744 VSS.n743 3.73383
R8220 VSS.n4505 VSS.n4504 3.73383
R8221 VSS.n2396 VSS.n2395 3.73383
R8222 VSS.n1981 VSS.n1702 3.73383
R8223 VSS.n3072 VSS.n1443 3.73383
R8224 VSS.n2727 VSS.n2622 3.73383
R8225 VSS.n3159 VSS.n1389 3.73383
R8226 VSS.n4446 VSS.n847 3.73383
R8227 VSS.n1342 VSS.n1341 3.73383
R8228 VSS.n1318 VSS.n901 3.73383
R8229 VSS.n53 VSS.n49 3.70885
R8230 VSS.n4064 VSS.n61 3.6913
R8231 VSS.n2394 VSS.n383 3.6029
R8232 VSS.n5445 VSS.n113 3.55606
R8233 VSS.n4832 VSS.n638 3.55606
R8234 VSS.n2361 VSS.n2067 3.55606
R8235 VSS.n2470 VSS.n1701 3.55606
R8236 VSS.n3056 VSS.n1456 3.55606
R8237 VSS.n328 VSS.n295 3.55606
R8238 VSS.n4199 VSS.n4198 3.55606
R8239 VSS.n1957 VSS.n1956 3.55606
R8240 VSS.n1436 VSS.n1435 3.55606
R8241 VSS.n5377 VSS.n239 3.55606
R8242 VSS.n2620 VSS.n2619 3.53424
R8243 VSS.n2924 VSS.n2922 3.53424
R8244 VSS.n1625 VSS.n1624 3.53424
R8245 VSS.n5222 VSS.n405 3.53424
R8246 VSS.n2174 VSS.n2173 3.53424
R8247 VSS.n1925 VSS.n393 3.53424
R8248 VSS.n2873 VSS.n2870 3.53424
R8249 VSS.n3228 VSS.n3225 3.53424
R8250 VSS.n3897 VSS.n947 3.53424
R8251 VSS.n3190 VSS.n3189 3.53424
R8252 VSS.n4472 VSS.n840 3.53424
R8253 VSS.n1386 VSS.n1385 3.53424
R8254 VSS.n1892 VSS.n1891 3.53424
R8255 VSS.n706 VSS.n705 3.53424
R8256 VSS.n4679 VSS.n672 3.53424
R8257 VSS.n3805 VSS.n3802 3.53424
R8258 VSS.n4402 VSS.n961 3.53424
R8259 VSS.n3283 VSS.n3282 3.53424
R8260 VSS.n4227 VSS.n4226 3.53424
R8261 VSS.n3308 VSS.n151 3.53424
R8262 VSS.n4014 VSS.n1128 3.33889
R8263 VSS.n2925 VSS.n2924 3.29866
R8264 VSS.n5223 VSS.n5222 3.29866
R8265 VSS.n5227 VSS.n393 3.29866
R8266 VSS.n3256 VSS.n3255 3.29866
R8267 VSS.n4407 VSS.n947 3.29866
R8268 VSS.n4550 VSS.n840 3.29866
R8269 VSS.n3221 VSS.n3216 3.29866
R8270 VSS.n5122 VSS.n501 3.29866
R8271 VSS.n4781 VSS.n672 3.29866
R8272 VSS.n4403 VSS.n4402 3.29866
R8273 VSS.n3833 VSS.n3832 3.29866
R8274 VSS.n5427 VSS.n151 3.29866
R8275 VSS.n3256 VSS.n1347 3.22013
R8276 VSS.n3221 VSS.n3178 3.22013
R8277 VSS.n5122 VSS.n500 3.22013
R8278 VSS.n3833 VSS.n3801 3.22013
R8279 VSS.n4408 VSS.n900 3.1416
R8280 VSS.n839 VSS.n838 3.1416
R8281 VSS.n4782 VSS.n670 3.1416
R8282 VSS.n959 VSS.n958 3.1416
R8283 VSS.n1235 VSS 3.10518
R8284 VSS.n1287 VSS 3.10518
R8285 VSS VSS.n4515 3.10518
R8286 VSS VSS.n4621 3.10518
R8287 VSS VSS.n5084 3.10518
R8288 VSS.n1268 VSS.n1241 2.83284
R8289 VSS.n3925 VSS.n3924 2.83284
R8290 VSS.n4504 VSS.n4503 2.83284
R8291 VSS.n743 VSS.n737 2.83284
R8292 VSS.n5073 VSS.n5072 2.83284
R8293 VSS.n4329 VSS.n1013 2.82084
R8294 VSS.n1517 VSS.n335 2.82084
R8295 VSS.n2534 VSS.n1557 2.82084
R8296 VSS.n2290 VSS.n2222 2.82084
R8297 VSS.n2117 VSS.n2116 2.82084
R8298 VSS.t101 VSS.t54 2.78249
R8299 VSS.n3743 VSS.t90 2.78249
R8300 VSS.n4006 VSS.n4005 2.78249
R8301 VSS.n1270 VSS.n1269 2.77837
R8302 VSS.n3923 VSS.n3922 2.77837
R8303 VSS.n4493 VSS.n4463 2.77837
R8304 VSS.n736 VSS.n718 2.77837
R8305 VSS.n4331 VSS.n4330 2.7666
R8306 VSS.n1520 VSS.n1519 2.7666
R8307 VSS.n2533 VSS.n2532 2.7666
R8308 VSS.n2291 VSS.n2154 2.7666
R8309 VSS.n15 VSS.n0 2.7544
R8310 VSS.n76 VSS.n71 2.73369
R8311 VSS.n3348 VSS.n3340 2.73369
R8312 VSS.n2732 VSS.n246 2.73369
R8313 VSS.n5196 VSS.n419 2.73369
R8314 VSS.n1952 VSS.n1916 2.73369
R8315 VSS.n4119 VSS.n28 2.73369
R8316 VSS.n5362 VSS.n304 2.73369
R8317 VSS.n5370 VSS.n294 2.73369
R8318 VSS.n1681 VSS.n1680 2.73369
R8319 VSS.n2465 VSS.n2001 2.73369
R8320 VSS.n1271 VSS.n1270 2.7239
R8321 VSS.n3922 VSS.n898 2.7239
R8322 VSS.n4493 VSS.n785 2.7239
R8323 VSS.n4656 VSS.n718 2.7239
R8324 VSS.n4102 VSS.n4067 2.71236
R8325 VSS.n4101 VSS.n4068 2.71236
R8326 VSS.n4077 VSS.n4074 2.71236
R8327 VSS.n4095 VSS.n4094 2.71236
R8328 VSS.n4091 VSS.n4078 2.71236
R8329 VSS.n4090 VSS.n4079 2.71236
R8330 VSS.n4084 VSS.n4083 2.71236
R8331 VSS.n4080 VSS.n1016 2.71236
R8332 VSS.n4323 VSS.n4322 2.71236
R8333 VSS.n4398 VSS.n4331 2.71236
R8334 VSS.n4337 VSS.n4336 2.71236
R8335 VSS.n4391 VSS.n4390 2.71236
R8336 VSS.n4365 VSS.n4338 2.71236
R8337 VSS.n4364 VSS.n4340 2.71236
R8338 VSS.n4359 VSS.n4358 2.71236
R8339 VSS.n4354 VSS.n4342 2.71236
R8340 VSS.n4353 VSS.n4346 2.71236
R8341 VSS.n4348 VSS.n4347 2.71236
R8342 VSS.n5294 VSS.n334 2.71236
R8343 VSS.n1521 VSS.n1520 2.71236
R8344 VSS.n2561 VSS.n1489 2.71236
R8345 VSS.n2560 VSS.n1490 2.71236
R8346 VSS.n1531 VSS.n1528 2.71236
R8347 VSS.n2554 VSS.n2553 2.71236
R8348 VSS.n2550 VSS.n1532 2.71236
R8349 VSS.n2549 VSS.n1533 2.71236
R8350 VSS.n1540 VSS.n1537 2.71236
R8351 VSS.n2543 VSS.n2542 2.71236
R8352 VSS.n2539 VSS.n1541 2.71236
R8353 VSS.n2532 VSS.n2531 2.71236
R8354 VSS.n1567 VSS.n1566 2.71236
R8355 VSS.n2523 VSS.n2522 2.71236
R8356 VSS.n2232 VSS.n1568 2.71236
R8357 VSS.n2237 VSS.n2236 2.71236
R8358 VSS.n2242 VSS.n2231 2.71236
R8359 VSS.n2243 VSS.n2229 2.71236
R8360 VSS.n2250 VSS.n2248 2.71236
R8361 VSS.n2249 VSS.n2226 2.71236
R8362 VSS.n2284 VSS.n2283 2.71236
R8363 VSS.n2294 VSS.n2154 2.71236
R8364 VSS.n2301 VSS.n2299 2.71236
R8365 VSS.n2300 VSS.n2128 2.71236
R8366 VSS.n2308 VSS.n2307 2.71236
R8367 VSS.n2130 VSS.n2129 2.71236
R8368 VSS.n2317 VSS.n2124 2.71236
R8369 VSS.n2316 VSS.n2122 2.71236
R8370 VSS.n2323 VSS.n2121 2.71236
R8371 VSS.n2325 VSS.n2324 2.71236
R8372 VSS.n2332 VSS.n2115 2.71236
R8373 VSS.n5064 VSS.n583 2.69529
R8374 VSS.n1178 VSS.n1177 2.65147
R8375 VSS.n5014 VSS.n609 2.61497
R8376 VSS.n3992 VSS.n3991 2.61497
R8377 VSS.n3956 VSS.n3955 2.61497
R8378 VSS.n4425 VSS.n4424 2.61497
R8379 VSS.n4604 VSS.n4603 2.61497
R8380 VSS.n4655 VSS.n734 2.61497
R8381 VSS.n4066 VSS.n4065 2.60389
R8382 VSS.n4397 VSS.n4332 2.60389
R8383 VSS.n1522 VSS.n1488 2.60389
R8384 VSS.n2529 VSS.n1562 2.60389
R8385 VSS.n2295 VSS.n2152 2.60389
R8386 VSS.n3337 VSS.n3335 2.59839
R8387 VSS.n5376 VSS.n241 2.59839
R8388 VSS.n1434 VSS.n416 2.59839
R8389 VSS.n1955 VSS.n1954 2.59839
R8390 VSS.n4990 VSS.n628 2.59839
R8391 VSS.n4254 VSS.n4253 2.59839
R8392 VSS.n5367 VSS.n5366 2.59839
R8393 VSS.n3055 VSS.n1458 2.59839
R8394 VSS.n2469 VSS.n1997 2.59839
R8395 VSS.n5256 VSS.n364 2.59839
R8396 VSS.n3993 VSS.n1215 2.58636
R8397 VSS.n5015 VSS.n608 2.58636
R8398 VSS.n5544 VSS.n28 2.45707
R8399 VSS.n5481 VSS.n71 2.45707
R8400 VSS.n5262 VSS.n360 2.45707
R8401 VSS.n4982 VSS.n4952 2.45707
R8402 VSS.n4009 VSS.n4008 2.38255
R8403 VSS.n3991 VSS.n3990 2.28816
R8404 VSS.n3955 VSS.n3954 2.28816
R8405 VSS.n4424 VSS.n892 2.28816
R8406 VSS.n4603 VSS.n779 2.28816
R8407 VSS.n734 VSS.n561 2.28816
R8408 VSS.n4067 VSS.n4066 2.27847
R8409 VSS.n4336 VSS.n4332 2.27847
R8410 VSS.n1489 VSS.n1488 2.27847
R8411 VSS.n1566 VSS.n1562 2.27847
R8412 VSS.n2299 VSS.n2152 2.27847
R8413 VSS.n1174 VSS.n1166 2.25323
R8414 VSS VSS.n1191 2.24506
R8415 VSS.t12 VSS.n5 2.22609
R8416 VSS.t43 VSS.t29 2.22609
R8417 VSS.n1137 VSS.t41 2.22609
R8418 VSS.n4102 VSS.n4101 2.16999
R8419 VSS.n4074 VSS.n4068 2.16999
R8420 VSS.n4095 VSS.n4077 2.16999
R8421 VSS.n4094 VSS.n4078 2.16999
R8422 VSS.n4091 VSS.n4090 2.16999
R8423 VSS.n4084 VSS.n4079 2.16999
R8424 VSS.n4083 VSS.n4080 2.16999
R8425 VSS.n4323 VSS.n1016 2.16999
R8426 VSS.n4322 VSS.n1017 2.16999
R8427 VSS.n4391 VSS.n4337 2.16999
R8428 VSS.n4390 VSS.n4338 2.16999
R8429 VSS.n4365 VSS.n4364 2.16999
R8430 VSS.n4359 VSS.n4340 2.16999
R8431 VSS.n4358 VSS.n4342 2.16999
R8432 VSS.n4354 VSS.n4353 2.16999
R8433 VSS.n4348 VSS.n4346 2.16999
R8434 VSS.n4347 VSS.n334 2.16999
R8435 VSS.n5294 VSS.n5293 2.16999
R8436 VSS.n2561 VSS.n2560 2.16999
R8437 VSS.n1528 VSS.n1490 2.16999
R8438 VSS.n2554 VSS.n1531 2.16999
R8439 VSS.n2553 VSS.n1532 2.16999
R8440 VSS.n2550 VSS.n2549 2.16999
R8441 VSS.n1537 VSS.n1533 2.16999
R8442 VSS.n2543 VSS.n1540 2.16999
R8443 VSS.n2542 VSS.n1541 2.16999
R8444 VSS.n2539 VSS.n2538 2.16999
R8445 VSS.n2523 VSS.n1567 2.16999
R8446 VSS.n2522 VSS.n1568 2.16999
R8447 VSS.n2236 VSS.n2232 2.16999
R8448 VSS.n2237 VSS.n2231 2.16999
R8449 VSS.n2243 VSS.n2242 2.16999
R8450 VSS.n2248 VSS.n2229 2.16999
R8451 VSS.n2250 VSS.n2249 2.16999
R8452 VSS.n2284 VSS.n2226 2.16999
R8453 VSS.n2283 VSS.n2227 2.16999
R8454 VSS.n2301 VSS.n2300 2.16999
R8455 VSS.n2308 VSS.n2128 2.16999
R8456 VSS.n2307 VSS.n2130 2.16999
R8457 VSS.n2129 VSS.n2124 2.16999
R8458 VSS.n2317 VSS.n2316 2.16999
R8459 VSS.n2122 VSS.n2121 2.16999
R8460 VSS.n2325 VSS.n2323 2.16999
R8461 VSS.n2324 VSS.n2115 2.16999
R8462 VSS.n2332 VSS.n2331 2.16999
R8463 VSS.n2869 VSS.n2621 2.12075
R8464 VSS.n403 VSS.n402 2.12075
R8465 VSS.n392 VSS.n391 2.12075
R8466 VSS.n5428 VSS.n149 2.12075
R8467 VSS.n3965 VSS.n1241 2.07029
R8468 VSS.n3926 VSS.n3925 2.07029
R8469 VSS.n4504 VSS.n4444 2.07029
R8470 VSS.n743 VSS.n741 2.07029
R8471 VSS.n5073 VSS.n581 2.07029
R8472 VSS.n1017 VSS.n1013 2.06152
R8473 VSS.n5293 VSS.n335 2.06152
R8474 VSS.n2538 VSS.n1557 2.06152
R8475 VSS.n2227 VSS.n2222 2.06152
R8476 VSS.n2331 VSS.n2117 2.06152
R8477 VSS.n2925 VSS.n2869 1.8459
R8478 VSS.n5223 VSS.n403 1.8459
R8479 VSS.n5227 VSS.n392 1.8459
R8480 VSS.n5428 VSS.n5427 1.8459
R8481 VSS.n5514 VSS.n45 1.80664
R8482 VSS.n4018 VSS.n4017 1.80664
R8483 VSS.n3749 VSS.n3711 1.77399
R8484 VSS.n5232 VSS.n381 1.76337
R8485 VSS.n1199 VSS.t54 1.67753
R8486 VSS.t29 VSS.n5485 1.6697
R8487 VSS.n3756 VSS.n3579 1.61978
R8488 VSS.n1172 VSS.n1171 1.607
R8489 VSS.n1179 VSS.n1178 1.5546
R8490 VSS.n4018 VSS.n1115 1.49252
R8491 VSS.n4881 VSS.n609 1.41667
R8492 VSS.n4775 VSS.n4774 1.41667
R8493 VSS.n3335 VSS.n113 1.40769
R8494 VSS.n5377 VSS.n5376 1.40769
R8495 VSS.n1435 VSS.n1434 1.40769
R8496 VSS.n1956 VSS.n1955 1.40769
R8497 VSS.n4832 VSS.n628 1.40769
R8498 VSS.n4254 VSS.n4199 1.40769
R8499 VSS.n5366 VSS.n295 1.40769
R8500 VSS.n3056 VSS.n3055 1.40769
R8501 VSS.n2470 VSS.n2469 1.40769
R8502 VSS.n2361 VSS.n364 1.40769
R8503 VSS.n3337 VSS.n3333 1.38063
R8504 VSS.n2897 VSS.n241 1.38063
R8505 VSS.n5197 VSS.n416 1.38063
R8506 VSS.n1954 VSS.n1953 1.38063
R8507 VSS.n4253 VSS.n4252 1.38063
R8508 VSS.n5367 VSS.n293 1.38063
R8509 VSS.n1613 VSS.n1458 1.38063
R8510 VSS.n2199 VSS.n1997 1.38063
R8511 VSS.n3340 VSS.n3333 1.35357
R8512 VSS.n2897 VSS.n246 1.35357
R8513 VSS.n5197 VSS.n5196 1.35357
R8514 VSS.n1953 VSS.n1952 1.35357
R8515 VSS.n4252 VSS.n304 1.35357
R8516 VSS.n5370 VSS.n293 1.35357
R8517 VSS.n1680 VSS.n1613 1.35357
R8518 VSS.n2199 VSS.n2001 1.35357
R8519 VSS.n4774 VSS.n594 1.30773
R8520 VSS.n4046 VSS.n76 1.29944
R8521 VSS.n3349 VSS.n3348 1.29944
R8522 VSS.n2733 VSS.n2732 1.29944
R8523 VSS.n440 VSS.n419 1.29944
R8524 VSS.n1916 VSS.n664 1.29944
R8525 VSS.n4120 VSS.n4119 1.29944
R8526 VSS.n5362 VSS.n5361 1.29944
R8527 VSS.n2578 VSS.n294 1.29944
R8528 VSS.n1681 VSS.n1575 1.29944
R8529 VSS.n2465 VSS.n2464 1.29944
R8530 VSS.n1270 VSS.n1267 1.29343
R8531 VSS.n4494 VSS.n4493 1.29343
R8532 VSS.n3922 VSS.n3921 1.29343
R8533 VSS.n4660 VSS.n718 1.29343
R8534 VSS.n1953 VSS.n1880 1.22878
R8535 VSS.n2200 VSS.n2199 1.22878
R8536 VSS.n1676 VSS.n1613 1.22878
R8537 VSS.n1494 VSS.n293 1.22878
R8538 VSS.n4252 VSS.n4224 1.22878
R8539 VSS.n2898 VSS.n2897 1.22878
R8540 VSS.n5198 VSS.n5197 1.22878
R8541 VSS.n3333 VSS.n3332 1.22878
R8542 VSS.n3506 VSS.n3505 1.14433
R8543 VSS.n2774 VSS.n2745 1.14433
R8544 VSS.n4409 VSS.n867 1.14433
R8545 VSS.n4551 VSS.n786 1.14433
R8546 VSS.n3177 VSS.n447 1.14433
R8547 VSS.n4802 VSS.n4801 1.14433
R8548 VSS.n4783 VSS.n538 1.14433
R8549 VSS.n3761 VSS.n3760 1.14433
R8550 VSS.n3425 VSS.n3421 1.14433
R8551 VSS.n4024 VSS.n4023 1.14433
R8552 VSS.n163 VSS.n148 1.13948
R8553 VSS.n2868 VSS.n2585 1.13948
R8554 VSS.n1742 VSS.n1723 1.13948
R8555 VSS.n2432 VSS.n2431 1.13948
R8556 VSS.n4141 VSS.n4138 1.13948
R8557 VSS.n4046 VSS.n4045 1.13708
R8558 VSS.n3349 VSS.n191 1.13708
R8559 VSS.n2735 VSS.n2733 1.13708
R8560 VSS.n440 VSS.n439 1.13708
R8561 VSS.n664 VSS.n658 1.13708
R8562 VSS.n4120 VSS.n1039 1.13708
R8563 VSS.n5361 VSS.n5360 1.13708
R8564 VSS.n2578 VSS.n1485 1.13708
R8565 VSS.n1577 VSS.n1575 1.13708
R8566 VSS.n2464 VSS.n2463 1.13708
R8567 VSS.n4015 VSS.t32 1.1133
R8568 VSS.n3368 VSS.n3367 1.08986
R8569 VSS.n3499 VSS.n3372 1.08986
R8570 VSS.n3412 VSS.n3411 1.08986
R8571 VSS.n3407 VSS.n3378 1.08986
R8572 VSS.n3380 VSS.n3379 1.08986
R8573 VSS.n3402 VSS.n3384 1.08986
R8574 VSS.n3396 VSS.n3395 1.08986
R8575 VSS.n3391 VSS.n3390 1.08986
R8576 VSS.n3840 VSS.n3839 1.08986
R8577 VSS.n2790 VSS.n2773 1.08986
R8578 VSS.n2770 VSS.n2747 1.08986
R8579 VSS.n2767 VSS.n2766 1.08986
R8580 VSS.n2754 VSS.n2749 1.08986
R8581 VSS.n2759 VSS.n2756 1.08986
R8582 VSS.n3146 VSS.n1411 1.08986
R8583 VSS.n1415 VSS.n1412 1.08986
R8584 VSS.n3153 VSS.n3152 1.08986
R8585 VSS.n3158 VSS.n3156 1.08986
R8586 VSS.n4536 VSS.n868 1.08986
R8587 VSS.n941 VSS.n906 1.08986
R8588 VSS.n909 VSS.n908 1.08986
R8589 VSS.n936 VSS.n910 1.08986
R8590 VSS.n933 VSS.n932 1.08986
R8591 VSS.n927 VSS.n918 1.08986
R8592 VSS.n922 VSS.n921 1.08986
R8593 VSS.n4544 VSS.n844 1.08986
R8594 VSS.n4445 VSS.n845 1.08986
R8595 VSS.n4586 VSS.n4585 1.08986
R8596 VSS.n4581 VSS.n794 1.08986
R8597 VSS.n798 VSS.n797 1.08986
R8598 VSS.n4576 VSS.n799 1.08986
R8599 VSS.n4573 VSS.n4572 1.08986
R8600 VSS.n4568 VSS.n809 1.08986
R8601 VSS.n813 VSS.n812 1.08986
R8602 VSS.n4563 VSS.n814 1.08986
R8603 VSS.n4560 VSS.n4559 1.08986
R8604 VSS.n5156 VSS.n448 1.08986
R8605 VSS.n5153 VSS.n5152 1.08986
R8606 VSS.n5130 VSS.n455 1.08986
R8607 VSS.n5146 VSS.n458 1.08986
R8608 VSS.n486 VSS.n459 1.08986
R8609 VSS.n5135 VSS.n467 1.08986
R8610 VSS.n5139 VSS.n468 1.08986
R8611 VSS.n495 VSS.n494 1.08986
R8612 VSS.n5127 VSS.n5126 1.08986
R8613 VSS.n5117 VSS.n510 1.08986
R8614 VSS.n515 VSS.n511 1.08986
R8615 VSS.n5111 VSS.n516 1.08986
R8616 VSS.n4850 VSS.n4846 1.08986
R8617 VSS.n4859 VSS.n4843 1.08986
R8618 VSS.n4864 VSS.n4863 1.08986
R8619 VSS.n4868 VSS.n4867 1.08986
R8620 VSS.n4873 VSS.n4872 1.08986
R8621 VSS.n5105 VSS.n539 1.08986
R8622 VSS.n4743 VSS.n4730 1.08986
R8623 VSS.n4745 VSS.n4728 1.08986
R8624 VSS.n4750 VSS.n4726 1.08986
R8625 VSS.n4753 VSS.n4727 1.08986
R8626 VSS.n4758 VSS.n4725 1.08986
R8627 VSS.n4761 VSS.n4724 1.08986
R8628 VSS.n4769 VSS.n4768 1.08986
R8629 VSS.n4776 VSS.n4692 1.08986
R8630 VSS.n3653 VSS.n3649 1.08986
R8631 VSS.n3657 VSS.n3616 1.08986
R8632 VSS.n3662 VSS.n3615 1.08986
R8633 VSS.n3666 VSS.n3614 1.08986
R8634 VSS.n3671 VSS.n3613 1.08986
R8635 VSS.n3675 VSS.n3612 1.08986
R8636 VSS.n3676 VSS.n3611 1.08986
R8637 VSS.n3681 VSS.n3589 1.08986
R8638 VSS.n3706 VSS.n3590 1.08986
R8639 VSS.n3477 VSS.n3423 1.08986
R8640 VSS.n3474 VSS.n3473 1.08986
R8641 VSS.n3451 VSS.n3448 1.08986
R8642 VSS.n3461 VSS.n3455 1.08986
R8643 VSS.n3465 VSS.n3457 1.08986
R8644 VSS.n3865 VSS.n1314 1.08986
R8645 VSS.n1316 VSS.n1315 1.08986
R8646 VSS.n3872 VSS.n3871 1.08986
R8647 VSS.n1306 VSS.n1305 1.08986
R8648 VSS.n3783 VSS.n3782 1.08986
R8649 VSS.n3793 VSS.n3527 1.08986
R8650 VSS.n3530 VSS.n3528 1.08986
R8651 VSS.n3788 VSS.n3532 1.08986
R8652 VSS.n3554 VSS.n3553 1.08986
R8653 VSS.n3574 VSS.n3573 1.08986
R8654 VSS.n3561 VSS.n3559 1.08986
R8655 VSS.n3567 VSS.n3565 1.08986
R8656 VSS.n3799 VSS.n3523 1.08986
R8657 VSS.n5422 VSS.n161 1.08525
R8658 VSS.n168 VSS.n162 1.08525
R8659 VSS.n5416 VSS.n169 1.08525
R8660 VSS.n2653 VSS.n2651 1.08525
R8661 VSS.n2657 VSS.n2655 1.08525
R8662 VSS.n2665 VSS.n2664 1.08525
R8663 VSS.n2669 VSS.n2668 1.08525
R8664 VSS.n2720 VSS.n2646 1.08525
R8665 VSS.n2726 VSS.n2639 1.08525
R8666 VSS.n2968 VSS.n2586 1.08525
R8667 VSS.n2964 VSS.n2963 1.08525
R8668 VSS.n2937 VSS.n2936 1.08525
R8669 VSS.n2957 VSS.n2932 1.08525
R8670 VSS.n2941 VSS.n2933 1.08525
R8671 VSS.n2951 VSS.n2943 1.08525
R8672 VSS.n3078 VSS.n1447 1.08525
R8673 VSS.n1449 VSS.n1448 1.08525
R8674 VSS.n3086 VSS.n3085 1.08525
R8675 VSS.n1766 VSS.n1721 1.08525
R8676 VSS.n1773 VSS.n1771 1.08525
R8677 VSS.n1780 VSS.n1779 1.08525
R8678 VSS.n1718 VSS.n1716 1.08525
R8679 VSS.n1786 VSS.n1717 1.08525
R8680 VSS.n1792 VSS.n1791 1.08525
R8681 VSS.n1800 VSS.n1799 1.08525
R8682 VSS.n1706 VSS.n1703 1.08525
R8683 VSS.n1977 VSS.n1705 1.08525
R8684 VSS.n2038 VSS.n2034 1.08525
R8685 VSS.n2420 VSS.n2042 1.08525
R8686 VSS.n2423 VSS.n2419 1.08525
R8687 VSS.n2415 VSS.n2044 1.08525
R8688 VSS.n2051 VSS.n2047 1.08525
R8689 VSS.n2405 VSS.n2055 1.08525
R8690 VSS.n2408 VSS.n2404 1.08525
R8691 VSS.n2400 VSS.n2057 1.08525
R8692 VSS.n2393 VSS.n2060 1.08525
R8693 VSS.n4150 VSS.n1061 1.08525
R8694 VSS.n4152 VSS.n1057 1.08525
R8695 VSS.n4156 VSS.n1058 1.08525
R8696 VSS.n1083 VSS.n1080 1.08525
R8697 VSS.n1088 VSS.n1078 1.08525
R8698 VSS.n1093 VSS.n1092 1.08525
R8699 VSS.n1073 VSS.n1069 1.08525
R8700 VSS.n1103 VSS.n1068 1.08525
R8701 VSS.n1100 VSS.n147 1.08525
R8702 VSS.n5470 VSS.n84 1.08295
R8703 VSS.n89 VSS.n85 1.08295
R8704 VSS.n5464 VSS.n90 1.08295
R8705 VSS.n126 VSS.n124 1.08295
R8706 VSS.n130 VSS.n128 1.08295
R8707 VSS.n135 VSS.n121 1.08295
R8708 VSS.n138 VSS.n118 1.08295
R8709 VSS.n5452 VSS.n5451 1.08295
R8710 VSS.n5459 VSS.n5458 1.08295
R8711 VSS.n5410 VSS.n192 1.08295
R8712 VSS.n5407 VSS.n5406 1.08295
R8713 VSS.n5402 VSS.n200 1.08295
R8714 VSS.n5398 VSS.n201 1.08295
R8715 VSS.n228 VSS.n223 1.08295
R8716 VSS.n5393 VSS.n5392 1.08295
R8717 VSS.n5388 VSS.n232 1.08295
R8718 VSS.n5384 VSS.n5382 1.08295
R8719 VSS.n5378 VSS.n236 1.08295
R8720 VSS.n2848 VSS.n2736 1.08295
R8721 VSS.n2845 VSS.n2844 1.08295
R8722 VSS.n2829 VSS.n2828 1.08295
R8723 VSS.n2838 VSS.n2818 1.08295
R8724 VSS.n2833 VSS.n2819 1.08295
R8725 VSS.n3111 VSS.n1429 1.08295
R8726 VSS.n1431 VSS.n1430 1.08295
R8727 VSS.n3120 VSS.n3119 1.08295
R8728 VSS.n1433 VSS.n1421 1.08295
R8729 VSS.n5186 VSS.n429 1.08295
R8730 VSS.n434 VSS.n430 1.08295
R8731 VSS.n5180 VSS.n435 1.08295
R8732 VSS.n1825 VSS.n1823 1.08295
R8733 VSS.n1829 VSS.n1827 1.08295
R8734 VSS.n1839 VSS.n1838 1.08295
R8735 VSS.n1817 VSS.n1816 1.08295
R8736 VSS.n1871 VSS.n1869 1.08295
R8737 VSS.n1877 VSS.n1810 1.08295
R8738 VSS.n4936 VSS.n662 1.08295
R8739 VSS.n4933 VSS.n4932 1.08295
R8740 VSS.n4928 VSS.n4825 1.08295
R8741 VSS.n4924 VSS.n4826 1.08295
R8742 VSS.n4920 VSS.n4919 1.08295
R8743 VSS.n4912 VSS.n4911 1.08295
R8744 VSS.n4904 VSS.n4903 1.08295
R8745 VSS.n4944 VSS.n635 1.08295
R8746 VSS.n4831 VSS.n636 1.08295
R8747 VSS.n4316 VSS.n1040 1.08295
R8748 VSS.n4280 VSS.n4267 1.08295
R8749 VSS.n4282 VSS.n4265 1.08295
R8750 VSS.n4287 VSS.n4263 1.08295
R8751 VSS.n4290 VSS.n4264 1.08295
R8752 VSS.n4295 VSS.n4262 1.08295
R8753 VSS.n4298 VSS.n4261 1.08295
R8754 VSS.n4304 VSS.n4303 1.08295
R8755 VSS.n4311 VSS.n4310 1.08295
R8756 VSS.n317 VSS.n307 1.08295
R8757 VSS.n5348 VSS.n311 1.08295
R8758 VSS.n5352 VSS.n312 1.08295
R8759 VSS.n5323 VSS.n5322 1.08295
R8760 VSS.n2683 VSS.n2681 1.08295
R8761 VSS.n2694 VSS.n2693 1.08295
R8762 VSS.n2687 VSS.n2677 1.08295
R8763 VSS.n5316 VSS.n323 1.08295
R8764 VSS.n326 VSS.n325 1.08295
R8765 VSS.n3041 VSS.n1486 1.08295
R8766 VSS.n3038 VSS.n3037 1.08295
R8767 VSS.n3009 VSS.n3008 1.08295
R8768 VSS.n3031 VSS.n2998 1.08295
R8769 VSS.n3000 VSS.n2999 1.08295
R8770 VSS.n3026 VSS.n3004 1.08295
R8771 VSS.n3022 VSS.n3021 1.08295
R8772 VSS.n3049 VSS.n1463 1.08295
R8773 VSS.n1464 VSS.n1457 1.08295
R8774 VSS.n2499 VSS.n1578 1.08295
R8775 VSS.n2496 VSS.n2495 1.08295
R8776 VSS.n2491 VSS.n1586 1.08295
R8777 VSS.n1591 VSS.n1587 1.08295
R8778 VSS.n2485 VSS.n1592 1.08295
R8779 VSS.n1692 VSS.n1691 1.08295
R8780 VSS.n2478 VSS.n2477 1.08295
R8781 VSS.n1697 VSS.n1696 1.08295
R8782 VSS.n2471 VSS.n1700 1.08295
R8783 VSS.n2459 VSS.n2006 1.08295
R8784 VSS.n2010 VSS.n2007 1.08295
R8785 VSS.n2453 VSS.n2011 1.08295
R8786 VSS.n2087 VSS.n2086 1.08295
R8787 VSS.n2092 VSS.n2091 1.08295
R8788 VSS.n2101 VSS.n2100 1.08295
R8789 VSS.n2106 VSS.n2105 1.08295
R8790 VSS.n2354 VSS.n2076 1.08295
R8791 VSS.n2360 VSS.n2068 1.08295
R8792 VSS.n3839 VSS.n1342 1.03539
R8793 VSS.n3159 VSS.n3158 1.03539
R8794 VSS.n4446 VSS.n4445 1.03539
R8795 VSS.n4559 VSS.n669 1.03539
R8796 VSS.n5126 VSS.n485 1.03539
R8797 VSS.n4881 VSS.n4880 1.03539
R8798 VSS.n4776 VSS.n4775 1.03539
R8799 VSS.n3706 VSS.n3705 1.03539
R8800 VSS.n1305 VSS.n901 1.03539
R8801 VSS.n3800 VSS.n3799 1.03539
R8802 VSS.n2727 VSS.n2726 1.03101
R8803 VSS.n3085 VSS.n1443 1.03101
R8804 VSS.n1705 VSS.n1702 1.03101
R8805 VSS.n2395 VSS.n2393 1.03101
R8806 VSS.n5429 VSS.n147 1.03101
R8807 VSS.n5458 VSS.n113 1.02883
R8808 VSS.n5378 VSS.n5377 1.02883
R8809 VSS.n1435 VSS.n1433 1.02883
R8810 VSS.n1956 VSS.n1877 1.02883
R8811 VSS.n4832 VSS.n4831 1.02883
R8812 VSS.n4310 VSS.n4199 1.02883
R8813 VSS.n325 VSS.n295 1.02883
R8814 VSS.n3056 VSS.n1457 1.02883
R8815 VSS.n2471 VSS.n2470 1.02883
R8816 VSS.n2361 VSS.n2360 1.02883
R8817 VSS.n3801 VSS.n3506 0.980926
R8818 VSS.n1347 VSS.n1342 0.980926
R8819 VSS.n2774 VSS.n1347 0.980926
R8820 VSS.n3178 VSS.n3159 0.980926
R8821 VSS.n4409 VSS.n4408 0.980926
R8822 VSS.n4446 VSS.n839 0.980926
R8823 VSS.n839 VSS.n786 0.980926
R8824 VSS.n4782 VSS.n669 0.980926
R8825 VSS.n3178 VSS.n3177 0.980926
R8826 VSS.n500 VSS.n485 0.980926
R8827 VSS.n4802 VSS.n500 0.980926
R8828 VSS.n4783 VSS.n4782 0.980926
R8829 VSS.n3761 VSS.n3579 0.980926
R8830 VSS.n3705 VSS.n959 0.980926
R8831 VSS.n3425 VSS.n959 0.980926
R8832 VSS.n4408 VSS.n901 0.980926
R8833 VSS.n4024 VSS.n1115 0.980926
R8834 VSS.n3801 VSS.n3800 0.980926
R8835 VSS.n5428 VSS.n148 0.976771
R8836 VSS.n2869 VSS.n2727 0.976771
R8837 VSS.n2869 VSS.n2868 0.976771
R8838 VSS.n1443 VSS.n403 0.976771
R8839 VSS.n1742 VSS.n403 0.976771
R8840 VSS.n1702 VSS.n392 0.976771
R8841 VSS.n2432 VSS.n392 0.976771
R8842 VSS.n2395 VSS.n2394 0.976771
R8843 VSS.n4138 VSS.n4064 0.976771
R8844 VSS.n5429 VSS.n5428 0.976771
R8845 VSS.n5539 VSS.n5538 0.975748
R8846 VSS.n5513 VSS.n46 0.975748
R8847 VSS.n5476 VSS.n5475 0.975748
R8848 VSS.n5231 VSS.n380 0.975748
R8849 VSS.n4954 VSS.n4951 0.975748
R8850 VSS.n615 VSS.n610 0.975748
R8851 VSS.n5041 VSS.n5040 0.975748
R8852 VSS.n5257 VSS.n363 0.975748
R8853 VSS.n3750 VSS.n3583 0.975748
R8854 VSS.n4016 VSS.n1125 0.975748
R8855 VSS.n3503 VSS.n3367 0.926457
R8856 VSS.n3500 VSS.n3499 0.926457
R8857 VSS.n3412 VSS.n3374 0.926457
R8858 VSS.n3378 VSS.n3377 0.926457
R8859 VSS.n3406 VSS.n3379 0.926457
R8860 VSS.n3396 VSS.n3386 0.926457
R8861 VSS.n3390 VSS.n3389 0.926457
R8862 VSS.n3840 VSS.n1324 0.926457
R8863 VSS.n2791 VSS.n2790 0.926457
R8864 VSS.n2771 VSS.n2770 0.926457
R8865 VSS.n2767 VSS.n2748 0.926457
R8866 VSS.n2764 VSS.n2749 0.926457
R8867 VSS.n2760 VSS.n2759 0.926457
R8868 VSS.n3145 VSS.n1415 0.926457
R8869 VSS.n3153 VSS.n1406 0.926457
R8870 VSS.n3156 VSS.n1405 0.926457
R8871 VSS.n4537 VSS.n4536 0.926457
R8872 VSS.n906 VSS.n905 0.926457
R8873 VSS.n940 VSS.n908 0.926457
R8874 VSS.n937 VSS.n936 0.926457
R8875 VSS.n933 VSS.n911 0.926457
R8876 VSS.n926 VSS.n921 0.926457
R8877 VSS.n923 VSS.n844 0.926457
R8878 VSS.n4543 VSS.n845 0.926457
R8879 VSS.n4586 VSS.n787 0.926457
R8880 VSS.n794 VSS.n790 0.926457
R8881 VSS.n4580 VSS.n797 0.926457
R8882 VSS.n4577 VSS.n4576 0.926457
R8883 VSS.n4573 VSS.n800 0.926457
R8884 VSS.n4567 VSS.n812 0.926457
R8885 VSS.n4564 VSS.n4563 0.926457
R8886 VSS.n4560 VSS.n833 0.926457
R8887 VSS.n5157 VSS.n5156 0.926457
R8888 VSS.n5153 VSS.n451 0.926457
R8889 VSS.n5130 VSS.n452 0.926457
R8890 VSS.n462 VSS.n458 0.926457
R8891 VSS.n5145 VSS.n459 0.926457
R8892 VSS.n5140 VSS.n5139 0.926457
R8893 VSS.n494 VSS.n493 0.926457
R8894 VSS.n5127 VSS.n484 0.926457
R8895 VSS.n4800 VSS.n510 0.926457
R8896 VSS.n5116 VSS.n511 0.926457
R8897 VSS.n5112 VSS.n5111 0.926457
R8898 VSS.n4846 VSS.n4845 0.926457
R8899 VSS.n4851 VSS.n4843 0.926457
R8900 VSS.n4867 VSS.n4841 0.926457
R8901 VSS.n4873 VSS.n4840 0.926457
R8902 VSS.n4876 VSS.n4839 0.926457
R8903 VSS.n5106 VSS.n5105 0.926457
R8904 VSS.n4730 VSS.n4729 0.926457
R8905 VSS.n4746 VSS.n4745 0.926457
R8906 VSS.n4750 VSS.n4749 0.926457
R8907 VSS.n4754 VSS.n4753 0.926457
R8908 VSS.n4762 VSS.n4761 0.926457
R8909 VSS.n4768 VSS.n4765 0.926457
R8910 VSS.n4770 VSS.n4692 0.926457
R8911 VSS VSS.n1234 0.926457
R8912 VSS VSS.n1285 0.926457
R8913 VSS.n4516 VSS 0.926457
R8914 VSS.n4622 VSS 0.926457
R8915 VSS.n5085 VSS 0.926457
R8916 VSS.n3649 VSS.n3580 0.926457
R8917 VSS.n3652 VSS.n3616 0.926457
R8918 VSS.n3658 VSS.n3615 0.926457
R8919 VSS.n3661 VSS.n3614 0.926457
R8920 VSS.n3667 VSS.n3613 0.926457
R8921 VSS.n3677 VSS.n3676 0.926457
R8922 VSS.n3681 VSS.n3680 0.926457
R8923 VSS.n3605 VSS.n3590 0.926457
R8924 VSS.n3478 VSS.n3477 0.926457
R8925 VSS.n3474 VSS.n3447 0.926457
R8926 VSS.n3471 VSS.n3448 0.926457
R8927 VSS.n3461 VSS.n3452 0.926457
R8928 VSS.n3466 VSS.n3465 0.926457
R8929 VSS.n3864 VSS.n1316 0.926457
R8930 VSS.n3872 VSS.n1308 0.926457
R8931 VSS.n1309 VSS.n1306 0.926457
R8932 VSS.n3783 VSS.n1116 0.926457
R8933 VSS.n3781 VSS.n3527 0.926457
R8934 VSS.n3792 VSS.n3528 0.926457
R8935 VSS.n3789 VSS.n3788 0.926457
R8936 VSS.n3555 VSS.n3554 0.926457
R8937 VSS.n3571 VSS.n3559 0.926457
R8938 VSS.n3568 VSS.n3567 0.926457
R8939 VSS.n3563 VSS.n3523 0.926457
R8940 VSS.n164 VSS.n161 0.922534
R8941 VSS.n5421 VSS.n162 0.922534
R8942 VSS.n5417 VSS.n5416 0.922534
R8943 VSS.n2651 VSS.n2650 0.922534
R8944 VSS.n2658 VSS.n2657 0.922534
R8945 VSS.n2668 VSS.n2648 0.922534
R8946 VSS.n2670 VSS.n2646 0.922534
R8947 VSS.n2719 VSS.n2639 0.922534
R8948 VSS.n2969 VSS.n2968 0.922534
R8949 VSS.n2964 VSS.n2589 0.922534
R8950 VSS.n2936 VSS.n2590 0.922534
R8951 VSS.n2938 VSS.n2932 0.922534
R8952 VSS.n2956 VSS.n2933 0.922534
R8953 VSS.n2942 VSS.n1447 0.922534
R8954 VSS.n3077 VSS.n1449 0.922534
R8955 VSS.n3086 VSS.n1442 0.922534
R8956 VSS.n1767 VSS.n1766 0.922534
R8957 VSS.n1771 VSS.n1770 0.922534
R8958 VSS.n1780 VSS.n1774 0.922534
R8959 VSS.n1777 VSS.n1718 0.922534
R8960 VSS.n1787 VSS.n1786 0.922534
R8961 VSS.n1800 VSS.n1708 0.922534
R8962 VSS.n1711 VSS.n1706 0.922534
R8963 VSS.n1978 VSS.n1977 0.922534
R8964 VSS.n2429 VSS.n2034 0.922534
R8965 VSS.n2420 VSS.n2036 0.922534
R8966 VSS.n2424 VSS.n2423 0.922534
R8967 VSS.n2044 VSS.n2043 0.922534
R8968 VSS.n2414 VSS.n2047 0.922534
R8969 VSS.n2409 VSS.n2408 0.922534
R8970 VSS.n2057 VSS.n2056 0.922534
R8971 VSS.n2399 VSS.n2060 0.922534
R8972 VSS.n4140 VSS.n1061 0.922534
R8973 VSS.n4152 VSS.n4151 0.922534
R8974 VSS.n4157 VSS.n4156 0.922534
R8975 VSS.n1080 VSS.n1079 0.922534
R8976 VSS.n1084 VSS.n1078 0.922534
R8977 VSS.n1077 VSS.n1069 0.922534
R8978 VSS.n1074 VSS.n1068 0.922534
R8979 VSS.n1102 VSS.n1100 0.922534
R8980 VSS.n4044 VSS.n84 0.920585
R8981 VSS.n5469 VSS.n85 0.920585
R8982 VSS.n5465 VSS.n5464 0.920585
R8983 VSS.n124 VSS.n123 0.920585
R8984 VSS.n131 VSS.n130 0.920585
R8985 VSS.n139 VSS.n138 0.920585
R8986 VSS.n5451 VSS.n5450 0.920585
R8987 VSS.n5459 VSS.n112 0.920585
R8988 VSS.n5411 VSS.n5410 0.920585
R8989 VSS.n5407 VSS.n195 0.920585
R8990 VSS.n200 VSS.n196 0.920585
R8991 VSS.n5401 VSS.n5398 0.920585
R8992 VSS.n224 VSS.n223 0.920585
R8993 VSS.n232 VSS.n220 0.920585
R8994 VSS.n5387 VSS.n5384 0.920585
R8995 VSS.n236 VSS.n233 0.920585
R8996 VSS.n2849 VSS.n2848 0.920585
R8997 VSS.n2845 VSS.n2811 0.920585
R8998 VSS.n2828 VSS.n2812 0.920585
R8999 VSS.n2830 VSS.n2818 0.920585
R9000 VSS.n2837 VSS.n2819 0.920585
R9001 VSS.n3110 VSS.n1431 0.920585
R9002 VSS.n3120 VSS.n1423 0.920585
R9003 VSS.n1424 VSS.n1421 0.920585
R9004 VSS.n438 VSS.n429 0.920585
R9005 VSS.n5185 VSS.n430 0.920585
R9006 VSS.n5181 VSS.n5180 0.920585
R9007 VSS.n1823 VSS.n1822 0.920585
R9008 VSS.n1827 VSS.n1826 0.920585
R9009 VSS.n1836 VSS.n1817 0.920585
R9010 VSS.n1869 VSS.n1815 0.920585
R9011 VSS.n1870 VSS.n1810 0.920585
R9012 VSS.n4937 VSS.n4936 0.920585
R9013 VSS.n4933 VSS.n4823 0.920585
R9014 VSS.n4825 VSS.n4824 0.920585
R9015 VSS.n4927 VSS.n4924 0.920585
R9016 VSS.n4920 VSS.n4829 0.920585
R9017 VSS.n4908 VSS.n4903 0.920585
R9018 VSS.n4905 VSS.n635 0.920585
R9019 VSS.n4943 VSS.n636 0.920585
R9020 VSS.n4317 VSS.n4316 0.920585
R9021 VSS.n4267 VSS.n4266 0.920585
R9022 VSS.n4283 VSS.n4282 0.920585
R9023 VSS.n4287 VSS.n4286 0.920585
R9024 VSS.n4291 VSS.n4290 0.920585
R9025 VSS.n4299 VSS.n4298 0.920585
R9026 VSS.n4303 VSS.n4302 0.920585
R9027 VSS.n4311 VSS.n4166 0.920585
R9028 VSS.n5358 VSS.n307 0.920585
R9029 VSS.n5348 VSS.n309 0.920585
R9030 VSS.n5353 VSS.n5352 0.920585
R9031 VSS.n5323 VSS.n314 0.920585
R9032 VSS.n2681 VSS.n315 0.920585
R9033 VSS.n2691 VSS.n2677 0.920585
R9034 VSS.n2688 VSS.n323 0.920585
R9035 VSS.n5315 VSS.n326 0.920585
R9036 VSS.n3042 VSS.n3041 0.920585
R9037 VSS.n3038 VSS.n2989 0.920585
R9038 VSS.n3009 VSS.n2990 0.920585
R9039 VSS.n3007 VSS.n2998 0.920585
R9040 VSS.n3030 VSS.n2999 0.920585
R9041 VSS.n3022 VSS.n3017 0.920585
R9042 VSS.n3020 VSS.n1463 0.920585
R9043 VSS.n3048 VSS.n1464 0.920585
R9044 VSS.n2500 VSS.n2499 0.920585
R9045 VSS.n2496 VSS.n1581 0.920585
R9046 VSS.n1586 VSS.n1582 0.920585
R9047 VSS.n2490 VSS.n1587 0.920585
R9048 VSS.n2486 VSS.n2485 0.920585
R9049 VSS.n2478 VSS.n1610 0.920585
R9050 VSS.n1696 VSS.n1611 0.920585
R9051 VSS.n2262 VSS.n1700 0.920585
R9052 VSS.n2006 VSS.n2004 0.920585
R9053 VSS.n2458 VSS.n2007 0.920585
R9054 VSS.n2454 VSS.n2453 0.920585
R9055 VSS.n2086 VSS.n2085 0.920585
R9056 VSS.n2093 VSS.n2092 0.920585
R9057 VSS.n2105 VSS.n2078 0.920585
R9058 VSS.n2107 VSS.n2076 0.920585
R9059 VSS.n2353 VSS.n2068 0.920585
R9060 VSS.n2621 VSS.n2620 0.903568
R9061 VSS.n1624 VSS.n402 0.903568
R9062 VSS.n2174 VSS.n391 0.903568
R9063 VSS.n2870 VSS.n1345 0.903568
R9064 VSS.n3225 VSS.n900 0.903568
R9065 VSS.n3189 VSS.n838 0.903568
R9066 VSS.n1386 VSS.n1355 0.903568
R9067 VSS.n1891 VSS.n498 0.903568
R9068 VSS.n705 VSS.n670 0.903568
R9069 VSS.n3802 VSS.n958 0.903568
R9070 VSS.n3282 VSS.n3263 0.903568
R9071 VSS.n4226 VSS.n149 0.903568
R9072 VSS.n3990 VSS.n1217 0.871989
R9073 VSS.n1223 VSS.n1222 0.871989
R9074 VSS.n3984 VSS.n3983 0.871989
R9075 VSS.n1226 VSS.n1224 0.871989
R9076 VSS.n3978 VSS.n1228 0.871989
R9077 VSS.n1236 VSS.n1235 0.871989
R9078 VSS.n3971 VSS.n3970 0.871989
R9079 VSS.n3966 VSS.n1237 0.871989
R9080 VSS.n3954 VSS.n3953 0.871989
R9081 VSS.n1277 VSS.n1275 0.871989
R9082 VSS.n3948 VSS.n1279 0.871989
R9083 VSS.n3947 VSS.n1280 0.871989
R9084 VSS.n3939 VSS.n3938 0.871989
R9085 VSS.n3933 VSS.n1287 0.871989
R9086 VSS.n3932 VSS.n1288 0.871989
R9087 VSS.n1296 VSS.n1295 0.871989
R9088 VSS.n4531 VSS.n892 0.871989
R9089 VSS.n4530 VSS.n893 0.871989
R9090 VSS.n4432 VSS.n4431 0.871989
R9091 VSS.n4524 VSS.n4523 0.871989
R9092 VSS.n4520 VSS.n4519 0.871989
R9093 VSS.n4515 VSS.n4434 0.871989
R9094 VSS.n4443 VSS.n4440 0.871989
R9095 VSS.n4509 VSS.n4508 0.871989
R9096 VSS.n4637 VSS.n779 0.871989
R9097 VSS.n4636 VSS.n780 0.871989
R9098 VSS.n4611 VSS.n4610 0.871989
R9099 VSS.n4630 VSS.n4629 0.871989
R9100 VSS.n4626 VSS.n4625 0.871989
R9101 VSS.n4621 VSS.n4616 0.871989
R9102 VSS.n4613 VSS.n740 0.871989
R9103 VSS.n4644 VSS.n4643 0.871989
R9104 VSS.n5100 VSS.n561 0.871989
R9105 VSS.n5099 VSS.n562 0.871989
R9106 VSS.n569 VSS.n568 0.871989
R9107 VSS.n5093 VSS.n5092 0.871989
R9108 VSS.n5089 VSS.n5088 0.871989
R9109 VSS.n5084 VSS.n571 0.871989
R9110 VSS.n580 VSS.n577 0.871989
R9111 VSS.n5078 VSS.n5077 0.871989
R9112 VSS.n4408 VSS.n4407 0.82504
R9113 VSS.n4550 VSS.n839 0.82504
R9114 VSS.n4782 VSS.n4781 0.82504
R9115 VSS.n4403 VSS.n959 0.82504
R9116 VSS.n5509 VSS.n5508 0.804553
R9117 VSS.n4007 VSS 0.786126
R9118 VSS.n4877 VSS.n4876 0.763053
R9119 VSS.n1347 VSS.n1345 0.746512
R9120 VSS.n3178 VSS.n1355 0.746512
R9121 VSS.n500 VSS.n498 0.746512
R9122 VSS.n3801 VSS.n3263 0.746512
R9123 VSS.n5505 VSS.n5504 0.686214
R9124 VSS.n5506 VSS.n5505 0.664786
R9125 VSS.n56 VSS.n55 0.664786
R9126 VSS.n1165 VSS.n1164 0.664786
R9127 VSS.n4011 VSS.n4010 0.664786
R9128 VSS.n30 VSS.n26 0.556899
R9129 VSS.n3977 VSS 0.545181
R9130 VSS VSS.n1283 0.545181
R9131 VSS VSS.n4433 0.545181
R9132 VSS VSS.n4612 0.545181
R9133 VSS VSS.n570 0.545181
R9134 VSS.n3403 VSS 0.463479
R9135 VSS VSS.n3402 0.463479
R9136 VSS.n2755 VSS 0.463479
R9137 VSS VSS.n1411 0.463479
R9138 VSS VSS.n917 0.463479
R9139 VSS.n918 VSS 0.463479
R9140 VSS VSS.n808 0.463479
R9141 VSS.n809 VSS 0.463479
R9142 VSS VSS.n465 0.463479
R9143 VSS.n5135 VSS 0.463479
R9144 VSS.n4858 VSS 0.463479
R9145 VSS.n4864 VSS 0.463479
R9146 VSS VSS.n4757 0.463479
R9147 VSS.n4758 VSS 0.463479
R9148 VSS.n3670 VSS 0.463479
R9149 VSS VSS.n3612 0.463479
R9150 VSS.n3456 VSS 0.463479
R9151 VSS VSS.n1314 0.463479
R9152 VSS VSS.n3558 0.463479
R9153 VSS.n3574 VSS 0.463479
R9154 VSS VSS.n2662 0.461517
R9155 VSS.n2665 VSS 0.461517
R9156 VSS.n2952 VSS 0.461517
R9157 VSS VSS.n2951 0.461517
R9158 VSS VSS.n1790 0.461517
R9159 VSS.n1791 VSS 0.461517
R9160 VSS VSS.n2049 0.461517
R9161 VSS.n2405 VSS 0.461517
R9162 VSS.n1087 VSS 0.461517
R9163 VSS.n1093 VSS 0.461517
R9164 VSS VSS.n134 0.460542
R9165 VSS.n135 VSS 0.460542
R9166 VSS.n227 VSS 0.460542
R9167 VSS.n5393 VSS 0.460542
R9168 VSS.n2834 VSS 0.460542
R9169 VSS VSS.n1429 0.460542
R9170 VSS.n1830 VSS 0.460542
R9171 VSS.n1839 VSS 0.460542
R9172 VSS.n4915 VSS 0.460542
R9173 VSS VSS.n4912 0.460542
R9174 VSS VSS.n4294 0.460542
R9175 VSS.n4295 VSS 0.460542
R9176 VSS.n2684 VSS 0.460542
R9177 VSS.n2694 VSS 0.460542
R9178 VSS.n3027 VSS 0.460542
R9179 VSS VSS.n3026 0.460542
R9180 VSS VSS.n1690 0.460542
R9181 VSS.n1691 VSS 0.460542
R9182 VSS VSS.n2097 0.460542
R9183 VSS.n2101 VSS 0.460542
R9184 VSS.n3505 VSS.n3503 0.436245
R9185 VSS.n3500 VSS.n3368 0.436245
R9186 VSS.n3374 VSS.n3372 0.436245
R9187 VSS.n3411 VSS.n3377 0.436245
R9188 VSS.n3407 VSS.n3406 0.436245
R9189 VSS.n3386 VSS.n3384 0.436245
R9190 VSS.n3395 VSS.n3389 0.436245
R9191 VSS.n3391 VSS.n1324 0.436245
R9192 VSS.n2791 VSS.n2745 0.436245
R9193 VSS.n2773 VSS.n2771 0.436245
R9194 VSS.n2748 VSS.n2747 0.436245
R9195 VSS.n2766 VSS.n2764 0.436245
R9196 VSS.n2760 VSS.n2754 0.436245
R9197 VSS.n3146 VSS.n3145 0.436245
R9198 VSS.n1412 VSS.n1406 0.436245
R9199 VSS.n3152 VSS.n1405 0.436245
R9200 VSS.n4537 VSS.n867 0.436245
R9201 VSS.n905 VSS.n868 0.436245
R9202 VSS.n941 VSS.n940 0.436245
R9203 VSS.n937 VSS.n909 0.436245
R9204 VSS.n911 VSS.n910 0.436245
R9205 VSS.n927 VSS.n926 0.436245
R9206 VSS.n923 VSS.n922 0.436245
R9207 VSS.n4544 VSS.n4543 0.436245
R9208 VSS.n4551 VSS.n787 0.436245
R9209 VSS.n4585 VSS.n790 0.436245
R9210 VSS.n4581 VSS.n4580 0.436245
R9211 VSS.n4577 VSS.n798 0.436245
R9212 VSS.n800 VSS.n799 0.436245
R9213 VSS.n4568 VSS.n4567 0.436245
R9214 VSS.n4564 VSS.n813 0.436245
R9215 VSS.n833 VSS.n814 0.436245
R9216 VSS.n5157 VSS.n447 0.436245
R9217 VSS.n451 VSS.n448 0.436245
R9218 VSS.n5152 VSS.n452 0.436245
R9219 VSS.n462 VSS.n455 0.436245
R9220 VSS.n5146 VSS.n5145 0.436245
R9221 VSS.n5140 VSS.n467 0.436245
R9222 VSS.n493 VSS.n468 0.436245
R9223 VSS.n495 VSS.n484 0.436245
R9224 VSS.n4801 VSS.n4800 0.436245
R9225 VSS.n5117 VSS.n5116 0.436245
R9226 VSS.n5112 VSS.n515 0.436245
R9227 VSS.n4845 VSS.n516 0.436245
R9228 VSS.n4851 VSS.n4850 0.436245
R9229 VSS.n4863 VSS.n4841 0.436245
R9230 VSS.n4868 VSS.n4840 0.436245
R9231 VSS.n4872 VSS.n4839 0.436245
R9232 VSS.n5106 VSS.n538 0.436245
R9233 VSS.n4729 VSS.n539 0.436245
R9234 VSS.n4746 VSS.n4743 0.436245
R9235 VSS.n4749 VSS.n4728 0.436245
R9236 VSS.n4754 VSS.n4726 0.436245
R9237 VSS.n4762 VSS.n4725 0.436245
R9238 VSS.n4765 VSS.n4724 0.436245
R9239 VSS.n4770 VSS.n4769 0.436245
R9240 VSS.n3760 VSS.n3580 0.436245
R9241 VSS.n3653 VSS.n3652 0.436245
R9242 VSS.n3658 VSS.n3657 0.436245
R9243 VSS.n3662 VSS.n3661 0.436245
R9244 VSS.n3667 VSS.n3666 0.436245
R9245 VSS.n3677 VSS.n3675 0.436245
R9246 VSS.n3680 VSS.n3611 0.436245
R9247 VSS.n3605 VSS.n3589 0.436245
R9248 VSS.n3478 VSS.n3421 0.436245
R9249 VSS.n3447 VSS.n3423 0.436245
R9250 VSS.n3473 VSS.n3471 0.436245
R9251 VSS.n3452 VSS.n3451 0.436245
R9252 VSS.n3466 VSS.n3455 0.436245
R9253 VSS.n3865 VSS.n3864 0.436245
R9254 VSS.n1315 VSS.n1308 0.436245
R9255 VSS.n3871 VSS.n1309 0.436245
R9256 VSS.n4023 VSS.n1116 0.436245
R9257 VSS.n3782 VSS.n3781 0.436245
R9258 VSS.n3793 VSS.n3792 0.436245
R9259 VSS.n3789 VSS.n3530 0.436245
R9260 VSS.n3555 VSS.n3532 0.436245
R9261 VSS.n3573 VSS.n3571 0.436245
R9262 VSS.n3568 VSS.n3561 0.436245
R9263 VSS.n3565 VSS.n3563 0.436245
R9264 VSS.n164 VSS.n163 0.434398
R9265 VSS.n5422 VSS.n5421 0.434398
R9266 VSS.n5417 VSS.n168 0.434398
R9267 VSS.n2650 VSS.n169 0.434398
R9268 VSS.n2658 VSS.n2653 0.434398
R9269 VSS.n2664 VSS.n2648 0.434398
R9270 VSS.n2670 VSS.n2669 0.434398
R9271 VSS.n2720 VSS.n2719 0.434398
R9272 VSS.n2969 VSS.n2585 0.434398
R9273 VSS.n2589 VSS.n2586 0.434398
R9274 VSS.n2963 VSS.n2590 0.434398
R9275 VSS.n2938 VSS.n2937 0.434398
R9276 VSS.n2957 VSS.n2956 0.434398
R9277 VSS.n2943 VSS.n2942 0.434398
R9278 VSS.n3078 VSS.n3077 0.434398
R9279 VSS.n1448 VSS.n1442 0.434398
R9280 VSS.n1767 VSS.n1723 0.434398
R9281 VSS.n1770 VSS.n1721 0.434398
R9282 VSS.n1774 VSS.n1773 0.434398
R9283 VSS.n1779 VSS.n1777 0.434398
R9284 VSS.n1787 VSS.n1716 0.434398
R9285 VSS.n1792 VSS.n1708 0.434398
R9286 VSS.n1799 VSS.n1711 0.434398
R9287 VSS.n1978 VSS.n1703 0.434398
R9288 VSS.n2431 VSS.n2429 0.434398
R9289 VSS.n2038 VSS.n2036 0.434398
R9290 VSS.n2424 VSS.n2042 0.434398
R9291 VSS.n2419 VSS.n2043 0.434398
R9292 VSS.n2415 VSS.n2414 0.434398
R9293 VSS.n2409 VSS.n2055 0.434398
R9294 VSS.n2404 VSS.n2056 0.434398
R9295 VSS.n2400 VSS.n2399 0.434398
R9296 VSS.n4141 VSS.n4140 0.434398
R9297 VSS.n4151 VSS.n4150 0.434398
R9298 VSS.n4157 VSS.n1057 0.434398
R9299 VSS.n1079 VSS.n1058 0.434398
R9300 VSS.n1084 VSS.n1083 0.434398
R9301 VSS.n1092 VSS.n1077 0.434398
R9302 VSS.n1074 VSS.n1073 0.434398
R9303 VSS.n1103 VSS.n1102 0.434398
R9304 VSS.n4045 VSS.n4044 0.433481
R9305 VSS.n5470 VSS.n5469 0.433481
R9306 VSS.n5465 VSS.n89 0.433481
R9307 VSS.n123 VSS.n90 0.433481
R9308 VSS.n131 VSS.n126 0.433481
R9309 VSS.n139 VSS.n121 0.433481
R9310 VSS.n5450 VSS.n118 0.433481
R9311 VSS.n5452 VSS.n112 0.433481
R9312 VSS.n5411 VSS.n191 0.433481
R9313 VSS.n195 VSS.n192 0.433481
R9314 VSS.n5406 VSS.n196 0.433481
R9315 VSS.n5402 VSS.n5401 0.433481
R9316 VSS.n224 VSS.n201 0.433481
R9317 VSS.n5392 VSS.n220 0.433481
R9318 VSS.n5388 VSS.n5387 0.433481
R9319 VSS.n5382 VSS.n233 0.433481
R9320 VSS.n2849 VSS.n2735 0.433481
R9321 VSS.n2811 VSS.n2736 0.433481
R9322 VSS.n2844 VSS.n2812 0.433481
R9323 VSS.n2830 VSS.n2829 0.433481
R9324 VSS.n2838 VSS.n2837 0.433481
R9325 VSS.n3111 VSS.n3110 0.433481
R9326 VSS.n1430 VSS.n1423 0.433481
R9327 VSS.n3119 VSS.n1424 0.433481
R9328 VSS.n439 VSS.n438 0.433481
R9329 VSS.n5186 VSS.n5185 0.433481
R9330 VSS.n5181 VSS.n434 0.433481
R9331 VSS.n1822 VSS.n435 0.433481
R9332 VSS.n1826 VSS.n1825 0.433481
R9333 VSS.n1838 VSS.n1836 0.433481
R9334 VSS.n1816 VSS.n1815 0.433481
R9335 VSS.n1871 VSS.n1870 0.433481
R9336 VSS.n4937 VSS.n658 0.433481
R9337 VSS.n4823 VSS.n662 0.433481
R9338 VSS.n4932 VSS.n4824 0.433481
R9339 VSS.n4928 VSS.n4927 0.433481
R9340 VSS.n4829 VSS.n4826 0.433481
R9341 VSS.n4911 VSS.n4908 0.433481
R9342 VSS.n4905 VSS.n4904 0.433481
R9343 VSS.n4944 VSS.n4943 0.433481
R9344 VSS.n4317 VSS.n1039 0.433481
R9345 VSS.n4266 VSS.n1040 0.433481
R9346 VSS.n4283 VSS.n4280 0.433481
R9347 VSS.n4286 VSS.n4265 0.433481
R9348 VSS.n4291 VSS.n4263 0.433481
R9349 VSS.n4299 VSS.n4262 0.433481
R9350 VSS.n4302 VSS.n4261 0.433481
R9351 VSS.n4304 VSS.n4166 0.433481
R9352 VSS.n5360 VSS.n5358 0.433481
R9353 VSS.n317 VSS.n309 0.433481
R9354 VSS.n5353 VSS.n311 0.433481
R9355 VSS.n314 VSS.n312 0.433481
R9356 VSS.n5322 VSS.n315 0.433481
R9357 VSS.n2693 VSS.n2691 0.433481
R9358 VSS.n2688 VSS.n2687 0.433481
R9359 VSS.n5316 VSS.n5315 0.433481
R9360 VSS.n3042 VSS.n1485 0.433481
R9361 VSS.n2989 VSS.n1486 0.433481
R9362 VSS.n3037 VSS.n2990 0.433481
R9363 VSS.n3008 VSS.n3007 0.433481
R9364 VSS.n3031 VSS.n3030 0.433481
R9365 VSS.n3017 VSS.n3004 0.433481
R9366 VSS.n3021 VSS.n3020 0.433481
R9367 VSS.n3049 VSS.n3048 0.433481
R9368 VSS.n2500 VSS.n1577 0.433481
R9369 VSS.n1581 VSS.n1578 0.433481
R9370 VSS.n2495 VSS.n1582 0.433481
R9371 VSS.n2491 VSS.n2490 0.433481
R9372 VSS.n2486 VSS.n1591 0.433481
R9373 VSS.n1692 VSS.n1610 0.433481
R9374 VSS.n2477 VSS.n1611 0.433481
R9375 VSS.n2262 VSS.n1697 0.433481
R9376 VSS.n2463 VSS.n2004 0.433481
R9377 VSS.n2459 VSS.n2458 0.433481
R9378 VSS.n2454 VSS.n2010 0.433481
R9379 VSS.n2085 VSS.n2011 0.433481
R9380 VSS.n2093 VSS.n2087 0.433481
R9381 VSS.n2100 VSS.n2078 0.433481
R9382 VSS.n2107 VSS.n2106 0.433481
R9383 VSS.n2354 VSS.n2353 0.433481
R9384 VSS.n4008 VSS.n4007 0.33298
R9385 VSS.n4880 VSS.n4877 0.327309
R9386 VSS.n1234 VSS 0.327309
R9387 VSS.n1285 VSS 0.327309
R9388 VSS.n4516 VSS 0.327309
R9389 VSS.n4622 VSS 0.327309
R9390 VSS.n5085 VSS 0.327309
R9391 VSS.n23 VSS.n15 0.320095
R9392 VSS.n19 VSS.n17 0.3165
R9393 VSS.n5506 VSS.n50 0.304763
R9394 VSS.n4010 VSS.n4009 0.285549
R9395 VSS.n5507 VSS.n5506 0.284166
R9396 VSS.n3380 VSS 0.27284
R9397 VSS.n2756 VSS 0.27284
R9398 VSS.n932 VSS 0.27284
R9399 VSS.n4572 VSS 0.27284
R9400 VSS.n486 VSS 0.27284
R9401 VSS.n4859 VSS 0.27284
R9402 VSS.n4727 VSS 0.27284
R9403 VSS.n3671 VSS 0.27284
R9404 VSS.n3457 VSS 0.27284
R9405 VSS.n3553 VSS 0.27284
R9406 VSS.n2655 VSS 0.271686
R9407 VSS VSS.n2941 0.271686
R9408 VSS.n1717 VSS 0.271686
R9409 VSS.n2051 VSS 0.271686
R9410 VSS.n1088 VSS 0.271686
R9411 VSS.n128 VSS 0.271113
R9412 VSS.n228 VSS 0.271113
R9413 VSS VSS.n2833 0.271113
R9414 VSS VSS.n1829 0.271113
R9415 VSS.n4919 VSS 0.271113
R9416 VSS.n4264 VSS 0.271113
R9417 VSS VSS.n2683 0.271113
R9418 VSS VSS.n3000 0.271113
R9419 VSS VSS.n1592 0.271113
R9420 VSS.n2091 VSS 0.271113
R9421 VSS.n24 VSS.n21 0.269191
R9422 VSS.n55 VSS.n54 0.26511
R9423 VSS.n5016 VSS.n5015 0.250777
R9424 VSS.n5566 VSS.n2 0.226306
R9425 VSS.n17 VSS.n2 0.1975
R9426 VSS.n1190 VSS.n48 0.18982
R9427 VSS.n1219 VSS.n48 0.18982
R9428 VSS.n1186 VSS.n1167 0.18982
R9429 VSS.n3403 VSS 0.163904
R9430 VSS VSS.n2755 0.163904
R9431 VSS.n917 VSS 0.163904
R9432 VSS.n808 VSS 0.163904
R9433 VSS VSS.n465 0.163904
R9434 VSS VSS.n4858 0.163904
R9435 VSS.n4757 VSS 0.163904
R9436 VSS VSS.n3670 0.163904
R9437 VSS VSS.n3456 0.163904
R9438 VSS.n3558 VSS 0.163904
R9439 VSS.n2662 VSS 0.163212
R9440 VSS.n2952 VSS 0.163212
R9441 VSS.n1790 VSS 0.163212
R9442 VSS VSS.n2049 0.163212
R9443 VSS VSS.n1087 0.163212
R9444 VSS.n134 VSS 0.162868
R9445 VSS VSS.n227 0.162868
R9446 VSS.n2834 VSS 0.162868
R9447 VSS.n1830 VSS 0.162868
R9448 VSS VSS.n4915 0.162868
R9449 VSS.n4294 VSS 0.162868
R9450 VSS.n2684 VSS 0.162868
R9451 VSS.n3027 VSS 0.162868
R9452 VSS.n1690 VSS 0.162868
R9453 VSS.n2097 VSS 0.162868
R9454 VSS.n21 VSS.n20 0.162714
R9455 VSS.n5510 VSS.n5509 0.148227
R9456 VSS.n5511 VSS.n5510 0.148227
R9457 VSS.n1189 VSS.n1188 0.148227
R9458 VSS.n1188 VSS.n1187 0.148227
R9459 VSS.n1177 VSS.n1176 0.0868708
R9460 VSS.n1176 VSS.n1175 0.0868708
R9461 VSS.n1175 VSS.n1174 0.0868708
R9462 VSS.n20 VSS.n19 0.0785
R9463 VSS.n23 VSS.n22 0.0665
R9464 VSS.n54 VSS.n53 0.0612955
R9465 VSS.n5015 VSS.n5014 0.0549681
R9466 VSS.n4990 VSS.n4952 0.0546226
R9467 VSS.n5256 VSS.n360 0.0546226
R9468 VSS.n2 VSS.n1 0.00533871
R9469 VSS.n24 VSS.n23 0.0035
R9470 w_18582_n15452.n0 w_18582_n15452.t28 433.272
R9471 w_18582_n15452.n0 w_18582_n15452.t15 433.272
R9472 w_18582_n15452.n0 w_18582_n15452.t27 433.149
R9473 w_18582_n15452.n0 w_18582_n15452.t20 433.149
R9474 w_18582_n15452.n0 w_18582_n15452.t24 433.149
R9475 w_18582_n15452.n0 w_18582_n15452.t21 433.149
R9476 w_18582_n15452.n0 w_18582_n15452.t17 433.149
R9477 w_18582_n15452.n0 w_18582_n15452.t14 433.149
R9478 w_18582_n15452.n0 w_18582_n15452.t26 433.149
R9479 w_18582_n15452.n0 w_18582_n15452.t23 433.149
R9480 w_18582_n15452.n0 w_18582_n15452.t18 433.149
R9481 w_18582_n15452.n0 w_18582_n15452.t16 433.149
R9482 w_18582_n15452.n0 w_18582_n15452.t13 433.149
R9483 w_18582_n15452.n0 w_18582_n15452.t25 433.149
R9484 w_18582_n15452.n0 w_18582_n15452.t22 433.149
R9485 w_18582_n15452.n0 w_18582_n15452.t19 433.149
R9486 w_18582_n15452.n1 w_18582_n15452.t10 228.546
R9487 w_18582_n15452.n1 w_18582_n15452.t12 228.215
R9488 w_18582_n15452.n1 w_18582_n15452.t6 228.215
R9489 w_18582_n15452.n1 w_18582_n15452.t8 228.215
R9490 w_18582_n15452.n3 w_18582_n15452.t0 216.696
R9491 w_18582_n15452.t5 w_18582_n15452.t11 173.161
R9492 w_18582_n15452.t7 w_18582_n15452.t9 173.161
R9493 w_18582_n15452.n5 w_18582_n15452.n4 154.19
R9494 w_18582_n15452.n6 w_18582_n15452.n5 152.655
R9495 w_18582_n15452.n2 w_18582_n15452.t5 86.5808
R9496 w_18582_n15452.n2 w_18582_n15452.t7 86.5808
R9497 w_18582_n15452.n1 w_18582_n15452.n2 48.0168
R9498 w_18582_n15452.n5 w_18582_n15452.n3 12.2118
R9499 w_18582_n15452.n0 w_18582_n15452.n1 7.57432
R9500 w_18582_n15452.n4 w_18582_n15452.t2 7.14175
R9501 w_18582_n15452.n4 w_18582_n15452.t3 7.14175
R9502 w_18582_n15452.t1 w_18582_n15452.n6 7.14175
R9503 w_18582_n15452.n6 w_18582_n15452.t4 7.14175
R9504 w_18582_n15452.n3 w_18582_n15452.n0 5.67084
R9505 MINUS.n4 MINUS.n2 167.306
R9506 MINUS.n4 MINUS.n3 167.091
R9507 MINUS.n12 MINUS.n11 83.5719
R9508 MINUS.n6 MINUS.t6 66.4617
R9509 MINUS.n5 MINUS.t7 66.1779
R9510 MINUS.n10 MINUS.t5 65.0304
R9511 MINUS.n13 MINUS.n12 64.9506
R9512 MINUS.n7 MINUS.t0 52.6863
R9513 MINUS.n3 MINUS.t3 5.7135
R9514 MINUS.n3 MINUS.t2 5.7135
R9515 MINUS.n2 MINUS.t1 5.7135
R9516 MINUS.n2 MINUS.t4 5.7135
R9517 MINUS.n8 MINUS.n4 3.41555
R9518 MINUS.n9 MINUS.n8 3.29465
R9519 MINUS.n11 MINUS.n10 1.56343
R9520 MINUS.n1 MINUS.n0 1.5505
R9521 MINUS.n13 MINUS.n1 1.33347
R9522 MINUS MINUS.n13 1.27403
R9523 MINUS.n11 MINUS.n0 0.77514
R9524 MINUS.n10 MINUS.n9 0.533273
R9525 MINUS.n7 MINUS.n6 0.5005
R9526 MINUS.n8 MINUS.n7 0.343415
R9527 MINUS MINUS.n0 0.314045
R9528 MINUS.n12 MINUS.t5 0.290206
R9529 MINUS.n5 MINUS 0.114798
R9530 MINUS.n6 MINUS.n5 0.083976
R9531 MINUS.n9 MINUS.n1 0.00690528
R9532 VDD.n28 VDD.t42 433.418
R9533 VDD.n9 VDD.t49 433.353
R9534 VDD.n41 VDD.t37 285.673
R9535 VDD.n29 VDD.t43 252.537
R9536 VDD.t40 VDD.n40 249.603
R9537 VDD.n8 VDD.t50 233.398
R9538 VDD.n3 VDD.t56 228.463
R9539 VDD.n0 VDD.t47 228.463
R9540 VDD.n3 VDD.t55 228.459
R9541 VDD.n0 VDD.t48 228.459
R9542 VDD.n2 VDD.t46 204.815
R9543 VDD.n5 VDD.t54 199.262
R9544 VDD.n33 VDD.t36 192.888
R9545 VDD.n38 VDD.t39 192.507
R9546 VDD.n9 VDD.t52 173.266
R9547 VDD.n28 VDD.t44 173.248
R9548 VDD.n11 VDD.n10 166.088
R9549 VDD.n13 VDD.n12 166.088
R9550 VDD.n15 VDD.n14 166.088
R9551 VDD.n17 VDD.n16 166.088
R9552 VDD.n19 VDD.n18 166.088
R9553 VDD.n21 VDD.n20 166.088
R9554 VDD.n23 VDD.n22 166.088
R9555 VDD.n25 VDD.n24 166.088
R9556 VDD.n27 VDD.n26 166.088
R9557 VDD.n32 VDD.t38 159.048
R9558 VDD.n39 VDD.t41 159.048
R9559 VDD.n35 VDD.n34 151.905
R9560 VDD.n37 VDD.n36 151.905
R9561 VDD.t57 VDD.t40 135.94
R9562 VDD.t0 VDD.t57 135.94
R9563 VDD.t59 VDD.t0 135.94
R9564 VDD.t34 VDD.t59 135.94
R9565 VDD.t37 VDD.t34 135.94
R9566 VDD.t28 VDD.t43 83.2968
R9567 VDD.t20 VDD.t28 83.2968
R9568 VDD.t14 VDD.t20 83.2968
R9569 VDD.t8 VDD.t14 83.2968
R9570 VDD.t32 VDD.t8 83.2968
R9571 VDD.t26 VDD.t32 83.2968
R9572 VDD.t22 VDD.t26 83.2968
R9573 VDD.t12 VDD.t22 83.2968
R9574 VDD.t6 VDD.t12 83.2968
R9575 VDD.t30 VDD.t6 83.2968
R9576 VDD.t24 VDD.t30 83.2968
R9577 VDD.t16 VDD.t24 83.2968
R9578 VDD.t10 VDD.t16 83.2968
R9579 VDD.t18 VDD.t10 83.2968
R9580 VDD.t4 VDD.t18 83.2968
R9581 VDD.t2 VDD.t4 83.2968
R9582 VDD.t50 VDD.t2 83.2968
R9583 VDD.n34 VDD.t60 7.14175
R9584 VDD.n34 VDD.t35 7.14175
R9585 VDD.n36 VDD.t58 7.14175
R9586 VDD.n36 VDD.t1 7.14175
R9587 VDD.n10 VDD.t3 5.7135
R9588 VDD.n10 VDD.t51 5.7135
R9589 VDD.n12 VDD.t19 5.7135
R9590 VDD.n12 VDD.t5 5.7135
R9591 VDD.n14 VDD.t17 5.7135
R9592 VDD.n14 VDD.t11 5.7135
R9593 VDD.n16 VDD.t31 5.7135
R9594 VDD.n16 VDD.t25 5.7135
R9595 VDD.n18 VDD.t13 5.7135
R9596 VDD.n18 VDD.t7 5.7135
R9597 VDD.n20 VDD.t27 5.7135
R9598 VDD.n20 VDD.t23 5.7135
R9599 VDD.n22 VDD.t9 5.7135
R9600 VDD.n22 VDD.t33 5.7135
R9601 VDD.n24 VDD.t21 5.7135
R9602 VDD.n24 VDD.t15 5.7135
R9603 VDD.n26 VDD.t44 5.7135
R9604 VDD.n26 VDD.t29 5.7135
R9605 VDD.n1 VDD.t45 4.93047
R9606 VDD.n4 VDD.t53 4.93036
R9607 VDD.n31 VDD.n30 2.29471
R9608 VDD VDD.n41 2.2075
R9609 VDD.n30 VDD.n29 2.15721
R9610 VDD.n40 VDD.n31 1.77198
R9611 VDD.n8 VDD.n7 1.69967
R9612 VDD.n6 VDD.n2 1.56377
R9613 VDD.n6 VDD.n5 0.782779
R9614 VDD.n7 VDD.n6 0.726584
R9615 VDD.n30 VDD.n7 0.290846
R9616 VDD.n37 VDD.n35 0.251473
R9617 VDD.n35 VDD.n33 0.205267
R9618 VDD.n38 VDD.n37 0.203807
R9619 VDD.n41 VDD.n32 0.153224
R9620 VDD.n27 VDD.n25 0.137178
R9621 VDD.n25 VDD.n23 0.137178
R9622 VDD.n23 VDD.n21 0.137178
R9623 VDD.n21 VDD.n19 0.137178
R9624 VDD.n19 VDD.n17 0.137178
R9625 VDD.n17 VDD.n15 0.137178
R9626 VDD.n15 VDD.n13 0.137178
R9627 VDD.n13 VDD.n11 0.137178
R9628 VDD.n40 VDD.n39 0.122095
R9629 VDD.n29 VDD.n28 0.12204
R9630 VDD.n9 VDD.n8 0.102565
R9631 VDD.n2 VDD.n1 0.0795521
R9632 VDD.n5 VDD.n4 0.0770473
R9633 VDD.n28 VDD.n27 0.0697042
R9634 VDD.n11 VDD.n9 0.067974
R9635 VDD.n39 VDD.n38 0.0481654
R9636 VDD.n33 VDD.n32 0.0467062
R9637 VDD VDD.n31 0.0272944
R9638 VDD.n4 VDD.n3 0.0185316
R9639 VDD.n1 VDD.n0 0.0184231
R9640 PLUS.n2 PLUS.n1 167.761
R9641 PLUS.n2 PLUS.n0 167.251
R9642 PLUS.n6 PLUS.t6 66.3341
R9643 PLUS.n8 PLUS.t7 66.1779
R9644 PLUS.n5 PLUS.t5 47.6794
R9645 PLUS.n3 PLUS.t0 47.4725
R9646 PLUS.n3 PLUS.n2 7.65247
R9647 PLUS.n1 PLUS.t3 5.7135
R9648 PLUS.n1 PLUS.t1 5.7135
R9649 PLUS.n0 PLUS.t2 5.7135
R9650 PLUS.n0 PLUS.t4 5.7135
R9651 PLUS.n7 PLUS.n4 4.78175
R9652 PLUS.n6 PLUS.n5 0.7505
R9653 PLUS.n8 PLUS.n7 0.21026
R9654 PLUS PLUS.n8 0.0801233
R9655 PLUS.n5 PLUS.n4 0.0790423
R9656 PLUS.n4 PLUS.n3 0.0547188
R9657 PLUS.n7 PLUS.n6 0.00178425
R9658 Gcm1 Gcm1.n1 213.453
R9659 Gcm1.n0 Gcm1.t7 192.851
R9660 Gcm1.n0 Gcm1.t6 192.851
R9661 Gcm1.n0 Gcm1.t2 192.475
R9662 Gcm1.n0 Gcm1.t0 192.475
R9663 Gcm1 Gcm1.n2 153.415
R9664 Gcm1.n2 Gcm1.t1 7.14175
R9665 Gcm1.n2 Gcm1.t3 7.14175
R9666 Gcm1 Gcm1.n0 5.50678
R9667 Gcm1.n1 Gcm1.t5 2.1755
R9668 Gcm1.n1 Gcm1.t4 2.1755
C0 a_12921_n6044# a_13253_n6644# 0.021022f
C1 a_14080_n6644# a_14246_n6044# 0.002572f
C2 a_13914_n6644# MINUS 0.00986f
C3 a_12589_n6644# PLUS 0.781424f
C4 a_19542_n12050# Gcm2 0.003537f
C5 VDD Gcm1 3.22615f
C6 VDD a_18606_n12050# 0.083842f
C7 a_13419_n6044# a_13914_n6644# 0.021323f
C8 a_19776_n11398# a_19308_n11398# 0.314775f
C9 a_13253_n6644# Sop 0.064431f
C10 a_19074_n12050# a_19308_n11398# 0.039502f
C11 a_13748_n6044# a_13914_n6644# 0.002479f
C12 a_12589_n6644# Gcm1 1.36e-19
C13 VDD a_12921_n6044# 0.023853f
C14 Vbgr PLUS 0.314462f
C15 a_14080_n6644# MINUS 0.089825f
C16 a_20010_n12050# a_20478_n12050# 0.314945f
C17 a_19308_n11398# Gcm2 0.03465f
C18 a_19776_n11398# a_20010_n12050# 0.038232f
C19 a_12589_n6644# a_12921_n6044# 0.021335f
C20 VDD Sop 0.029404f
C21 a_13087_n6644# MINUS 9.64e-20
C22 a_18840_n11398# XQ2[0|0].Emitter 8.03e-20
C23 a_13748_n6044# a_14080_n6644# 0.030096f
C24 VDD a_20478_n12050# 0.037731f
C25 a_13087_n6644# a_13419_n6044# 0.023472f
C26 VDD a_19776_n11398# 0.010539f
C27 a_12589_n6644# Sop 0.046808f
C28 a_20010_n12050# Gcm2 0.003343f
C29 VDD a_19074_n12050# 0.069535f
C30 VDD a_14246_n6044# 0.024218f
C31 a_13253_n6644# MINUS 0.00225f
C32 a_20244_n11398# a_19308_n11398# 3.64e-19
C33 PLUS Gcm1 0.857443f
C34 a_18606_n12050# PLUS 3.55e-19
C35 VDD Gcm2 1.60517f
C36 a_13253_n6644# a_13419_n6044# 0.008457f
C37 Vbgr a_20478_n12050# 0.04087f
C38 a_13253_n6644# a_13748_n6044# 0.023309f
C39 PLUS a_12921_n6044# 6.94e-19
C40 Vbgr a_19776_n11398# 4.33e-19
C41 VDD MINUS 2.53996f
C42 a_20010_n12050# a_20244_n11398# 0.039502f
C43 a_12755_n6044# a_13087_n6644# 0.030145f
C44 VDD a_13419_n6044# 0.030679f
C45 PLUS Sop 1.85175f
C46 VDD a_20244_n11398# 0.003996f
C47 VDD a_13748_n6044# 0.0148f
C48 Vbgr Gcm2 0.448781f
C49 a_20478_n12050# PLUS 2.58e-20
C50 a_19776_n11398# PLUS 0.002819f
C51 Gcm1 Sop 0.231375f
C52 a_19074_n12050# PLUS 4.12e-19
C53 Vbgr MINUS 0.870973f
C54 VDD XQ2[0|0].Emitter 0.16357f
C55 PLUS Gcm2 1.75721f
C56 a_12921_n6044# Sop 0.004563f
C57 VDD a_12755_n6044# 0.015049f
C58 a_18606_n12050# a_19074_n12050# 0.314564f
C59 Vbgr a_20244_n11398# 0.311719f
C60 a_13914_n6644# a_14080_n6644# 1.14572f
C61 PLUS MINUS 2.43119f
C62 a_12589_n6644# a_12755_n6044# 0.002355f
C63 a_18606_n12050# Gcm2 0.003522f
C64 a_13087_n6644# a_13914_n6644# 0.001343f
C65 PLUS a_13419_n6044# 2.08e-19
C66 a_18840_n11398# a_19308_n11398# 0.315392f
C67 Vbgr XQ2[0|0].Emitter 1.3e-19
C68 a_20244_n11398# PLUS 0.001875f
C69 Gcm1 MINUS 0.008743f
C70 Sop a_14246_n6044# 0.004293f
C71 a_12921_n6044# MINUS 6.48e-19
C72 a_13087_n6644# a_14080_n6644# 0.018599f
C73 a_13253_n6644# a_13914_n6644# 0.345538f
C74 a_19542_n12050# a_19308_n11398# 0.037557f
C75 Sop Gcm2 0.082758f
C76 PLUS XQ2[0|0].Emitter 0.223212f
C77 a_12921_n6044# a_13419_n6044# 0.355059f
C78 a_20478_n12050# Gcm2 0.003693f
C79 a_12755_n6044# PLUS 0.042938f
C80 a_19776_n11398# Gcm2 0.035089f
C81 Sop MINUS 1.99061f
C82 VDD a_18840_n11398# 0.022772f
C83 a_12921_n6044# a_13748_n6044# 1.29e-19
C84 a_19074_n12050# Gcm2 0.003576f
C85 VDD a_13914_n6644# 0.002202f
C86 a_19542_n12050# a_20010_n12050# 0.322063f
C87 a_13253_n6644# a_14080_n6644# 0.002946f
C88 a_13419_n6044# Sop 0.002172f
C89 Sop a_13748_n6044# 0.001245f
C90 a_12589_n6644# a_13914_n6644# 2.28e-19
C91 a_13087_n6644# a_13253_n6644# 0.921413f
C92 VDD a_19542_n12050# 0.070449f
C93 a_14246_n6044# MINUS 0.800786f
C94 a_20244_n11398# a_20478_n12050# 0.037563f
C95 a_19776_n11398# a_20244_n11398# 0.319832f
C96 VDD a_14080_n6644# 0.002932f
C97 a_12755_n6044# a_12921_n6044# 1.12551f
C98 Gcm2 MINUS 0.291314f
C99 a_13419_n6044# a_14246_n6044# 0.022788f
C100 a_13748_n6044# a_14246_n6044# 0.310596f
C101 VDD a_13087_n6644# 0.003097f
C102 a_12589_n6644# a_14080_n6644# 9.41e-22
C103 a_12755_n6044# Sop 3.93e-19
C104 a_20244_n11398# Gcm2 0.034686f
C105 VDD a_19308_n11398# 0.015546f
C106 a_12589_n6644# a_13087_n6644# 0.310844f
C107 a_13419_n6044# MINUS 0.003315f
C108 a_18840_n11398# PLUS 0.001491f
C109 a_13748_n6044# MINUS 0.040846f
C110 PLUS a_13914_n6644# 3.91e-19
C111 VDD a_13253_n6644# 0.002332f
C112 a_12755_n6044# a_14246_n6044# 3.01e-21
C113 VDD a_20010_n12050# 0.04598f
C114 a_13419_n6044# a_13748_n6044# 0.907295f
C115 a_18606_n12050# a_18840_n11398# 0.040276f
C116 a_12589_n6644# a_13253_n6644# 0.018593f
C117 a_19542_n12050# PLUS 4.28e-19
C118 XQ2[0|0].Emitter MINUS 4.53925f
C119 PLUS a_14080_n6644# 4.25e-20
C120 a_12755_n6044# MINUS 2.69e-19
C121 VDD a_12589_n6644# 0.002604f
C122 PLUS a_13087_n6644# 0.050677f
C123 a_12755_n6044# a_13419_n6044# 2.72e-19
C124 a_12755_n6044# a_13748_n6044# 0.018296f
C125 a_19308_n11398# PLUS 0.002747f
C126 Sop a_13914_n6644# 0.047735f
C127 VDD Vbgr 3.1251f
C128 PLUS a_13253_n6644# 0.005963f
C129 a_18840_n11398# a_19074_n12050# 0.037513f
C130 a_20010_n12050# PLUS 4.23e-19
C131 a_12921_n6044# a_13087_n6644# 0.002485f
C132 a_13914_n6644# a_14246_n6044# 0.021312f
C133 Sop a_14080_n6644# 0.011869f
C134 a_18840_n11398# Gcm2 0.034668f
C135 a_19542_n12050# a_19776_n11398# 0.039394f
C136 a_19542_n12050# a_19074_n12050# 0.315843f
C137 VDD PLUS 1.83264f
C138 a_13087_n6644# Sop 0.015632f
C139 Vbgr VSS 11.107247f
C140 VDD VSS 71.22097f
C141 a_20478_n12050# VSS 0.779933f
C142 a_20244_n11398# VSS 0.484218f
C143 a_20010_n12050# VSS 0.454007f
C144 a_19776_n11398# VSS 0.486416f
C145 a_19542_n12050# VSS 0.455174f
C146 a_19308_n11398# VSS 0.482581f
C147 a_19074_n12050# VSS 0.455714f
C148 a_18840_n11398# VSS 0.797756f
C149 a_18606_n12050# VSS 0.82397f
C150 XQ2[0|0].Emitter VSS 77.7933f
C151 Gcm2 VSS 3.40518f
C152 Sop VSS 5.80295f
C153 Gcm1 VSS 5.17281f
C154 MINUS VSS 7.397131f
C155 a_14246_n6044# VSS 0.89872f
C156 a_14080_n6644# VSS 0.754105f
C157 a_13914_n6644# VSS 0.512978f
C158 a_13748_n6044# VSS 0.637512f
C159 a_13419_n6044# VSS 0.797684f
C160 a_13253_n6644# VSS 0.71881f
C161 a_13087_n6644# VSS 0.602106f
C162 a_12921_n6044# VSS 0.567362f
C163 PLUS VSS 8.099231f
C164 a_12755_n6044# VSS 0.82331f
C165 a_12589_n6644# VSS 0.840352f
C166 Gcm1.n0 VSS 0.343643f
C167 Gcm1.t5 VSS 0.033806f
C168 Gcm1.t4 VSS 0.033806f
C169 Gcm1.n1 VSS 0.124907f
C170 Gcm1.t6 VSS 0.209367f
C171 Gcm1.t0 VSS 0.209207f
C172 Gcm1.t7 VSS 0.209367f
C173 Gcm1.t2 VSS 0.209207f
C174 Gcm1.t1 VSS 0.016903f
C175 Gcm1.t3 VSS 0.016903f
C176 Gcm1.n2 VSS 0.051633f
C177 PLUS.t2 VSS 0.006085f
C178 PLUS.t4 VSS 0.006085f
C179 PLUS.n0 VSS 0.019597f
C180 PLUS.t3 VSS 0.006085f
C181 PLUS.t1 VSS 0.006085f
C182 PLUS.n1 VSS 0.020001f
C183 PLUS.n2 VSS 0.511452f
C184 PLUS.t0 VSS 0.006494f
C185 PLUS.n3 VSS 0.336283f
C186 PLUS.n4 VSS 0.004602f
C187 PLUS.t6 VSS 0.438261f
C188 PLUS.t5 VSS 0.012875f
C189 PLUS.n5 VSS 0.122319f
C190 PLUS.n6 VSS 0.224294f
C191 PLUS.n7 VSS 0.031042f
C192 PLUS.t7 VSS 0.437785f
C193 PLUS.n8 VSS 0.173035f
C194 VDD.t45 VSS 0.360925f
C195 VDD.t48 VSS 0.006364f
C196 VDD.t47 VSS 0.006371f
C197 VDD.n0 VSS 0.533581f
C198 VDD.n1 VSS 0.128505f
C199 VDD.t46 VSS 0.605104f
C200 VDD.n2 VSS 0.724421f
C201 VDD.t54 VSS 0.597127f
C202 VDD.t56 VSS 0.006371f
C203 VDD.t55 VSS 0.006364f
C204 VDD.n3 VSS 0.533416f
C205 VDD.t53 VSS 0.360922f
C206 VDD.n4 VSS 0.125622f
C207 VDD.n5 VSS 0.500691f
C208 VDD.n6 VSS 0.86046f
C209 VDD.n7 VSS 0.298752f
C210 VDD.t43 VSS 0.238343f
C211 VDD.t42 VSS 0.051428f
C212 VDD.t44 VSS 0.051708f
C213 VDD.t49 VSS 0.051425f
C214 VDD.t52 VSS 0.043175f
C215 VDD.t28 VSS 0.167489f
C216 VDD.t20 VSS 0.167489f
C217 VDD.t14 VSS 0.167489f
C218 VDD.t8 VSS 0.167489f
C219 VDD.t32 VSS 0.167489f
C220 VDD.t26 VSS 0.167489f
C221 VDD.t22 VSS 0.167489f
C222 VDD.t12 VSS 0.167489f
C223 VDD.t6 VSS 0.167489f
C224 VDD.t30 VSS 0.167489f
C225 VDD.t24 VSS 0.167489f
C226 VDD.t16 VSS 0.167489f
C227 VDD.t10 VSS 0.167489f
C228 VDD.t18 VSS 0.167489f
C229 VDD.t4 VSS 0.167489f
C230 VDD.t2 VSS 0.167489f
C231 VDD.t50 VSS 0.327687f
C232 VDD.n8 VSS 0.26236f
C233 VDD.n9 VSS 0.088975f
C234 VDD.t3 VSS 0.00853f
C235 VDD.t51 VSS 0.00853f
C236 VDD.n10 VSS 0.027125f
C237 VDD.n11 VSS 0.049461f
C238 VDD.t19 VSS 0.00853f
C239 VDD.t5 VSS 0.00853f
C240 VDD.n12 VSS 0.027125f
C241 VDD.n13 VSS 0.063061f
C242 VDD.t17 VSS 0.00853f
C243 VDD.t11 VSS 0.00853f
C244 VDD.n14 VSS 0.027125f
C245 VDD.n15 VSS 0.063061f
C246 VDD.t31 VSS 0.00853f
C247 VDD.t25 VSS 0.00853f
C248 VDD.n16 VSS 0.027125f
C249 VDD.n17 VSS 0.063061f
C250 VDD.t13 VSS 0.00853f
C251 VDD.t7 VSS 0.00853f
C252 VDD.n18 VSS 0.027125f
C253 VDD.n19 VSS 0.063061f
C254 VDD.t27 VSS 0.00853f
C255 VDD.t23 VSS 0.00853f
C256 VDD.n20 VSS 0.027125f
C257 VDD.n21 VSS 0.063061f
C258 VDD.t9 VSS 0.00853f
C259 VDD.t33 VSS 0.00853f
C260 VDD.n22 VSS 0.027125f
C261 VDD.n23 VSS 0.063061f
C262 VDD.t21 VSS 0.00853f
C263 VDD.t15 VSS 0.00853f
C264 VDD.n24 VSS 0.027125f
C265 VDD.n25 VSS 0.063061f
C266 VDD.t29 VSS 0.00853f
C267 VDD.n26 VSS 0.027125f
C268 VDD.n27 VSS 0.0498f
C269 VDD.n28 VSS 0.093377f
C270 VDD.n29 VSS 0.136962f
C271 VDD.n30 VSS 1.24521f
C272 VDD.n31 VSS 0.993935f
C273 VDD.t38 VSS 0.033077f
C274 VDD.n32 VSS 0.041297f
C275 VDD.t39 VSS 0.084464f
C276 VDD.t36 VSS 0.084535f
C277 VDD.n33 VSS 0.075363f
C278 VDD.t60 VSS 0.006824f
C279 VDD.t35 VSS 0.006824f
C280 VDD.n34 VSS 0.020663f
C281 VDD.n35 VSS 0.079948f
C282 VDD.t58 VSS 0.006824f
C283 VDD.t1 VSS 0.006824f
C284 VDD.n36 VSS 0.020663f
C285 VDD.n37 VSS 0.079722f
C286 VDD.n38 VSS 0.07817f
C287 VDD.t41 VSS 0.033077f
C288 VDD.n39 VSS 0.036686f
C289 VDD.n40 VSS 0.438443f
C290 VDD.t40 VSS 0.418088f
C291 VDD.t57 VSS 0.273647f
C292 VDD.t0 VSS 0.273647f
C293 VDD.t59 VSS 0.273647f
C294 VDD.t34 VSS 0.273647f
C295 VDD.t37 VSS 0.448071f
C296 VDD.n41 VSS 0.556863f
C297 MINUS.n0 VSS 0.033171f
C298 MINUS.n1 VSS 0.480467f
C299 MINUS.t5 VSS 0.187676f
C300 MINUS.t1 VSS 0.023493f
C301 MINUS.t4 VSS 0.023493f
C302 MINUS.n2 VSS 0.075664f
C303 MINUS.t3 VSS 0.023493f
C304 MINUS.t2 VSS 0.023493f
C305 MINUS.n3 VSS 0.075679f
C306 MINUS.n4 VSS 1.4278f
C307 MINUS.t0 VSS 0.095737f
C308 MINUS.t6 VSS 1.69384f
C309 MINUS.t7 VSS 1.6902f
C310 MINUS.n5 VSS 0.617226f
C311 MINUS.n6 VSS 1.05159f
C312 MINUS.n7 VSS 0.779794f
C313 MINUS.n8 VSS 2.13651f
C314 MINUS.n9 VSS 1.18396f
C315 MINUS.n10 VSS 0.338979f
C316 MINUS.n11 VSS 0.085725f
C317 MINUS.n12 VSS 0.18589f
C318 MINUS.n13 VSS 0.276912f
C319 w_18582_n15452.t0 VSS 0.234962f
C320 w_18582_n15452.n0 VSS 3.48367f
C321 w_18582_n15452.n1 VSS 1.66094f
C322 w_18582_n15452.t4 VSS 0.021075f
C323 w_18582_n15452.t10 VSS 0.019545f
C324 w_18582_n15452.t8 VSS 0.019358f
C325 w_18582_n15452.t11 VSS 2.33369f
C326 w_18582_n15452.t5 VSS 1.42107f
C327 w_18582_n15452.t9 VSS 2.33369f
C328 w_18582_n15452.t7 VSS 1.42107f
C329 w_18582_n15452.n2 VSS 1.35891f
C330 w_18582_n15452.t6 VSS 0.019358f
C331 w_18582_n15452.t12 VSS 0.019358f
C332 w_18582_n15452.t15 VSS 0.158817f
C333 w_18582_n15452.t19 VSS 0.158794f
C334 w_18582_n15452.t22 VSS 0.158794f
C335 w_18582_n15452.t25 VSS 0.158794f
C336 w_18582_n15452.t13 VSS 0.158794f
C337 w_18582_n15452.t16 VSS 0.158794f
C338 w_18582_n15452.t18 VSS 0.158794f
C339 w_18582_n15452.t23 VSS 0.158794f
C340 w_18582_n15452.t26 VSS 0.158794f
C341 w_18582_n15452.t28 VSS 0.158817f
C342 w_18582_n15452.t27 VSS 0.158794f
C343 w_18582_n15452.t20 VSS 0.158794f
C344 w_18582_n15452.t24 VSS 0.158794f
C345 w_18582_n15452.t21 VSS 0.158794f
C346 w_18582_n15452.t17 VSS 0.158794f
C347 w_18582_n15452.t14 VSS 0.158794f
C348 w_18582_n15452.n3 VSS 1.23464f
C349 w_18582_n15452.t2 VSS 0.021075f
C350 w_18582_n15452.t3 VSS 0.021075f
C351 w_18582_n15452.n4 VSS 0.065747f
C352 w_18582_n15452.n5 VSS 0.884901f
C353 w_18582_n15452.n6 VSS 0.064031f
C354 w_18582_n15452.t1 VSS 0.021075f
C355 Vbgr.n0 VSS 0.005092f
C356 Vbgr.t2 VSS 0.022859f
C357 Vbgr.t1 VSS 0.022859f
C358 Vbgr.n1 VSS 0.072764f
C359 Vbgr.t0 VSS 0.022859f
C360 Vbgr.t3 VSS 0.022859f
C361 Vbgr.n2 VSS 0.07276f
C362 Vbgr.n3 VSS 0.461053f
C363 Vbgr.t4 VSS 0.037727f
C364 Vbgr.n4 VSS 0.048693f
C365 Vbgr.n5 VSS 0.186946f
C366 Vbgr.n6 VSS 0.040078f
C367 Vbgr.t6 VSS 0.978804f
C368 Vbgr.t7 VSS 0.965972f
C369 Vbgr.n7 VSS 2.31888f
C370 Vbgr.t8 VSS 0.965972f
C371 Vbgr.n8 VSS 1.17689f
C372 Vbgr.t5 VSS 0.965972f
C373 Vbgr.n9 VSS 1.7344f
C374 Vbgr.n10 VSS 0.336824f
C375 Vbgr.n11 VSS 0.008885f
.ends

